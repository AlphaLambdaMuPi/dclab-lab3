// Core.v

// Generated using ACDS version 15.1 185

`timescale 1 ps / 1 ps
module Core (
		inout  wire        audio_and_video_config_external_interface_SDAT,  // audio_and_video_config_external_interface.SDAT
		output wire        audio_and_video_config_external_interface_SCLK,  //                                          .SCLK
		input  wire        audio_external_interface_ADCDAT,                 //                  audio_external_interface.ADCDAT
		input  wire        audio_external_interface_ADCLRCK,                //                                          .ADCLRCK
		input  wire        audio_external_interface_BCLK,                   //                                          .BCLK
		output wire        audio_external_interface_DACDAT,                 //                                          .DACDAT
		input  wire        audio_external_interface_DACLRCK,                //                                          .DACLRCK
		input  wire        clk_clk,                                         //                                       clk.clk
		input  wire        clk_0_clk,                                       //                                     clk_0.clk
		output wire        clock_bridge_out_clk_clk,                        //                      clock_bridge_out_clk.clk
		input  wire        pio_touch_external_connection_export,            //             pio_touch_external_connection.export
		input  wire        reset_reset_n,                                   //                                     reset.reset_n
		input  wire        reset_0_reset_n,                                 //                                   reset_0.reset_n
		output wire [12:0] sdram_controller_wire_addr,                      //                     sdram_controller_wire.addr
		output wire [1:0]  sdram_controller_wire_ba,                        //                                          .ba
		output wire        sdram_controller_wire_cas_n,                     //                                          .cas_n
		output wire        sdram_controller_wire_cke,                       //                                          .cke
		output wire        sdram_controller_wire_cs_n,                      //                                          .cs_n
		inout  wire [31:0] sdram_controller_wire_dq,                        //                                          .dq
		output wire [3:0]  sdram_controller_wire_dqm,                       //                                          .dqm
		output wire        sdram_controller_wire_ras_n,                     //                                          .ras_n
		output wire        sdram_controller_wire_we_n,                      //                                          .we_n
		input  wire        spi_touch_external_MISO,                         //                        spi_touch_external.MISO
		output wire        spi_touch_external_MOSI,                         //                                          .MOSI
		output wire        spi_touch_external_SCLK,                         //                                          .SCLK
		output wire        spi_touch_external_SS_n,                         //                                          .SS_n
		inout  wire [15:0] sram_external_interface_DQ,                      //                   sram_external_interface.DQ
		output wire [19:0] sram_external_interface_ADDR,                    //                                          .ADDR
		output wire        sram_external_interface_LB_N,                    //                                          .LB_N
		output wire        sram_external_interface_UB_N,                    //                                          .UB_N
		output wire        sram_external_interface_CE_N,                    //                                          .CE_N
		output wire        sram_external_interface_OE_N,                    //                                          .OE_N
		output wire        sram_external_interface_WE_N,                    //                                          .WE_N
		output wire        sys_sdram_pll_sdram_clk_clk,                     //                   sys_sdram_pll_sdram_clk.clk
		output wire        video_vga_controller_external_interface_CLK,     //   video_vga_controller_external_interface.CLK
		output wire        video_vga_controller_external_interface_HS,      //                                          .HS
		output wire        video_vga_controller_external_interface_VS,      //                                          .VS
		output wire        video_vga_controller_external_interface_BLANK,   //                                          .BLANK
		output wire        video_vga_controller_external_interface_SYNC,    //                                          .SYNC
		output wire        video_vga_controller_external_interface_DATA_EN, //                                          .DATA_EN
		output wire [7:0]  video_vga_controller_external_interface_R,       //                                          .R
		output wire [7:0]  video_vga_controller_external_interface_G,       //                                          .G
		output wire [7:0]  video_vga_controller_external_interface_B        //                                          .B
	);

	wire         video_dual_clock_buffer_avalon_dc_buffer_source_valid;                       // video_dual_clock_buffer:stream_out_valid -> video_vga_controller:valid
	wire  [29:0] video_dual_clock_buffer_avalon_dc_buffer_source_data;                        // video_dual_clock_buffer:stream_out_data -> video_vga_controller:data
	wire         video_dual_clock_buffer_avalon_dc_buffer_source_ready;                       // video_vga_controller:ready -> video_dual_clock_buffer:stream_out_ready
	wire         video_dual_clock_buffer_avalon_dc_buffer_source_startofpacket;               // video_dual_clock_buffer:stream_out_startofpacket -> video_vga_controller:startofpacket
	wire         video_dual_clock_buffer_avalon_dc_buffer_source_endofpacket;                 // video_dual_clock_buffer:stream_out_endofpacket -> video_vga_controller:endofpacket
	wire         video_pixel_buffer_dma_avalon_pixel_source_valid;                            // video_pixel_buffer_dma:stream_valid -> video_rgb_resampler_0:stream_in_valid
	wire  [15:0] video_pixel_buffer_dma_avalon_pixel_source_data;                             // video_pixel_buffer_dma:stream_data -> video_rgb_resampler_0:stream_in_data
	wire         video_pixel_buffer_dma_avalon_pixel_source_ready;                            // video_rgb_resampler_0:stream_in_ready -> video_pixel_buffer_dma:stream_ready
	wire         video_pixel_buffer_dma_avalon_pixel_source_startofpacket;                    // video_pixel_buffer_dma:stream_startofpacket -> video_rgb_resampler_0:stream_in_startofpacket
	wire         video_pixel_buffer_dma_avalon_pixel_source_endofpacket;                      // video_pixel_buffer_dma:stream_endofpacket -> video_rgb_resampler_0:stream_in_endofpacket
	wire         video_rgb_resampler_0_avalon_rgb_source_valid;                               // video_rgb_resampler_0:stream_out_valid -> video_dual_clock_buffer:stream_in_valid
	wire  [29:0] video_rgb_resampler_0_avalon_rgb_source_data;                                // video_rgb_resampler_0:stream_out_data -> video_dual_clock_buffer:stream_in_data
	wire         video_rgb_resampler_0_avalon_rgb_source_ready;                               // video_dual_clock_buffer:stream_in_ready -> video_rgb_resampler_0:stream_out_ready
	wire         video_rgb_resampler_0_avalon_rgb_source_startofpacket;                       // video_rgb_resampler_0:stream_out_startofpacket -> video_dual_clock_buffer:stream_in_startofpacket
	wire         video_rgb_resampler_0_avalon_rgb_source_endofpacket;                         // video_rgb_resampler_0:stream_out_endofpacket -> video_dual_clock_buffer:stream_in_endofpacket
	wire         video_pll_lcd_clk_clk;                                                       // video_pll:lcd_clk_clk -> [rst_controller_006:clk, rst_controller_007:clk, video_dual_clock_buffer:clk_stream_out, video_vga_controller:clk]
	wire         sys_sdram_pll_sys_clk_clk;                                                   // sys_sdram_pll:sys_clk_clk -> [irq_mapper:clk, irq_synchronizer:sender_clk, jtag_uart:clk, mm_interconnect_0:sys_sdram_pll_sys_clk_clk, nios2_cpu:clk, onchip_memory2:clk, pio_touch:clk, rst_controller_002:clk, rst_controller_004:clk, rst_controller_005:clk, sdram_controller:clk, spi_touch:clk, sram:clk, sysid_qsys:clock, timer:clk, video_dual_clock_buffer:clk_stream_in, video_pixel_buffer_dma:clk, video_rgb_resampler_0:clk]
	wire         video_pixel_buffer_dma_avalon_pixel_dma_master_waitrequest;                  // mm_interconnect_0:video_pixel_buffer_dma_avalon_pixel_dma_master_waitrequest -> video_pixel_buffer_dma:master_waitrequest
	wire  [15:0] video_pixel_buffer_dma_avalon_pixel_dma_master_readdata;                     // mm_interconnect_0:video_pixel_buffer_dma_avalon_pixel_dma_master_readdata -> video_pixel_buffer_dma:master_readdata
	wire  [31:0] video_pixel_buffer_dma_avalon_pixel_dma_master_address;                      // video_pixel_buffer_dma:master_address -> mm_interconnect_0:video_pixel_buffer_dma_avalon_pixel_dma_master_address
	wire         video_pixel_buffer_dma_avalon_pixel_dma_master_read;                         // video_pixel_buffer_dma:master_read -> mm_interconnect_0:video_pixel_buffer_dma_avalon_pixel_dma_master_read
	wire         video_pixel_buffer_dma_avalon_pixel_dma_master_readdatavalid;                // mm_interconnect_0:video_pixel_buffer_dma_avalon_pixel_dma_master_readdatavalid -> video_pixel_buffer_dma:master_readdatavalid
	wire         video_pixel_buffer_dma_avalon_pixel_dma_master_lock;                         // video_pixel_buffer_dma:master_arbiterlock -> mm_interconnect_0:video_pixel_buffer_dma_avalon_pixel_dma_master_lock
	wire  [31:0] nios2_cpu_data_master_readdata;                                              // mm_interconnect_0:nios2_cpu_data_master_readdata -> nios2_cpu:d_readdata
	wire         nios2_cpu_data_master_waitrequest;                                           // mm_interconnect_0:nios2_cpu_data_master_waitrequest -> nios2_cpu:d_waitrequest
	wire         nios2_cpu_data_master_debugaccess;                                           // nios2_cpu:debug_mem_slave_debugaccess_to_roms -> mm_interconnect_0:nios2_cpu_data_master_debugaccess
	wire  [28:0] nios2_cpu_data_master_address;                                               // nios2_cpu:d_address -> mm_interconnect_0:nios2_cpu_data_master_address
	wire   [3:0] nios2_cpu_data_master_byteenable;                                            // nios2_cpu:d_byteenable -> mm_interconnect_0:nios2_cpu_data_master_byteenable
	wire         nios2_cpu_data_master_read;                                                  // nios2_cpu:d_read -> mm_interconnect_0:nios2_cpu_data_master_read
	wire         nios2_cpu_data_master_readdatavalid;                                         // mm_interconnect_0:nios2_cpu_data_master_readdatavalid -> nios2_cpu:d_readdatavalid
	wire         nios2_cpu_data_master_write;                                                 // nios2_cpu:d_write -> mm_interconnect_0:nios2_cpu_data_master_write
	wire  [31:0] nios2_cpu_data_master_writedata;                                             // nios2_cpu:d_writedata -> mm_interconnect_0:nios2_cpu_data_master_writedata
	wire  [31:0] nios2_cpu_instruction_master_readdata;                                       // mm_interconnect_0:nios2_cpu_instruction_master_readdata -> nios2_cpu:i_readdata
	wire         nios2_cpu_instruction_master_waitrequest;                                    // mm_interconnect_0:nios2_cpu_instruction_master_waitrequest -> nios2_cpu:i_waitrequest
	wire  [28:0] nios2_cpu_instruction_master_address;                                        // nios2_cpu:i_address -> mm_interconnect_0:nios2_cpu_instruction_master_address
	wire         nios2_cpu_instruction_master_read;                                           // nios2_cpu:i_read -> mm_interconnect_0:nios2_cpu_instruction_master_read
	wire         nios2_cpu_instruction_master_readdatavalid;                                  // mm_interconnect_0:nios2_cpu_instruction_master_readdatavalid -> nios2_cpu:i_readdatavalid
	wire  [15:0] mm_interconnect_0_sram_avalon_sram_slave_readdata;                           // sram:readdata -> mm_interconnect_0:sram_avalon_sram_slave_readdata
	wire  [19:0] mm_interconnect_0_sram_avalon_sram_slave_address;                            // mm_interconnect_0:sram_avalon_sram_slave_address -> sram:address
	wire         mm_interconnect_0_sram_avalon_sram_slave_read;                               // mm_interconnect_0:sram_avalon_sram_slave_read -> sram:read
	wire   [1:0] mm_interconnect_0_sram_avalon_sram_slave_byteenable;                         // mm_interconnect_0:sram_avalon_sram_slave_byteenable -> sram:byteenable
	wire         mm_interconnect_0_sram_avalon_sram_slave_readdatavalid;                      // sram:readdatavalid -> mm_interconnect_0:sram_avalon_sram_slave_readdatavalid
	wire         mm_interconnect_0_sram_avalon_sram_slave_write;                              // mm_interconnect_0:sram_avalon_sram_slave_write -> sram:write
	wire  [15:0] mm_interconnect_0_sram_avalon_sram_slave_writedata;                          // mm_interconnect_0:sram_avalon_sram_slave_writedata -> sram:writedata
	wire         mm_interconnect_0_audio_avalon_audio_slave_chipselect;                       // mm_interconnect_0:audio_avalon_audio_slave_chipselect -> audio:chipselect
	wire  [31:0] mm_interconnect_0_audio_avalon_audio_slave_readdata;                         // audio:readdata -> mm_interconnect_0:audio_avalon_audio_slave_readdata
	wire   [1:0] mm_interconnect_0_audio_avalon_audio_slave_address;                          // mm_interconnect_0:audio_avalon_audio_slave_address -> audio:address
	wire         mm_interconnect_0_audio_avalon_audio_slave_read;                             // mm_interconnect_0:audio_avalon_audio_slave_read -> audio:read
	wire         mm_interconnect_0_audio_avalon_audio_slave_write;                            // mm_interconnect_0:audio_avalon_audio_slave_write -> audio:write
	wire  [31:0] mm_interconnect_0_audio_avalon_audio_slave_writedata;                        // mm_interconnect_0:audio_avalon_audio_slave_writedata -> audio:writedata
	wire  [31:0] mm_interconnect_0_audio_and_video_config_avalon_av_config_slave_readdata;    // audio_and_video_config:readdata -> mm_interconnect_0:audio_and_video_config_avalon_av_config_slave_readdata
	wire         mm_interconnect_0_audio_and_video_config_avalon_av_config_slave_waitrequest; // audio_and_video_config:waitrequest -> mm_interconnect_0:audio_and_video_config_avalon_av_config_slave_waitrequest
	wire   [1:0] mm_interconnect_0_audio_and_video_config_avalon_av_config_slave_address;     // mm_interconnect_0:audio_and_video_config_avalon_av_config_slave_address -> audio_and_video_config:address
	wire         mm_interconnect_0_audio_and_video_config_avalon_av_config_slave_read;        // mm_interconnect_0:audio_and_video_config_avalon_av_config_slave_read -> audio_and_video_config:read
	wire   [3:0] mm_interconnect_0_audio_and_video_config_avalon_av_config_slave_byteenable;  // mm_interconnect_0:audio_and_video_config_avalon_av_config_slave_byteenable -> audio_and_video_config:byteenable
	wire         mm_interconnect_0_audio_and_video_config_avalon_av_config_slave_write;       // mm_interconnect_0:audio_and_video_config_avalon_av_config_slave_write -> audio_and_video_config:write
	wire  [31:0] mm_interconnect_0_audio_and_video_config_avalon_av_config_slave_writedata;   // mm_interconnect_0:audio_and_video_config_avalon_av_config_slave_writedata -> audio_and_video_config:writedata
	wire  [31:0] mm_interconnect_0_video_pixel_buffer_dma_avalon_control_slave_readdata;      // video_pixel_buffer_dma:slave_readdata -> mm_interconnect_0:video_pixel_buffer_dma_avalon_control_slave_readdata
	wire   [1:0] mm_interconnect_0_video_pixel_buffer_dma_avalon_control_slave_address;       // mm_interconnect_0:video_pixel_buffer_dma_avalon_control_slave_address -> video_pixel_buffer_dma:slave_address
	wire         mm_interconnect_0_video_pixel_buffer_dma_avalon_control_slave_read;          // mm_interconnect_0:video_pixel_buffer_dma_avalon_control_slave_read -> video_pixel_buffer_dma:slave_read
	wire   [3:0] mm_interconnect_0_video_pixel_buffer_dma_avalon_control_slave_byteenable;    // mm_interconnect_0:video_pixel_buffer_dma_avalon_control_slave_byteenable -> video_pixel_buffer_dma:slave_byteenable
	wire         mm_interconnect_0_video_pixel_buffer_dma_avalon_control_slave_write;         // mm_interconnect_0:video_pixel_buffer_dma_avalon_control_slave_write -> video_pixel_buffer_dma:slave_write
	wire  [31:0] mm_interconnect_0_video_pixel_buffer_dma_avalon_control_slave_writedata;     // mm_interconnect_0:video_pixel_buffer_dma_avalon_control_slave_writedata -> video_pixel_buffer_dma:slave_writedata
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect;                    // mm_interconnect_0:jtag_uart_avalon_jtag_slave_chipselect -> jtag_uart:av_chipselect
	wire  [31:0] mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata;                      // jtag_uart:av_readdata -> mm_interconnect_0:jtag_uart_avalon_jtag_slave_readdata
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest;                   // jtag_uart:av_waitrequest -> mm_interconnect_0:jtag_uart_avalon_jtag_slave_waitrequest
	wire   [0:0] mm_interconnect_0_jtag_uart_avalon_jtag_slave_address;                       // mm_interconnect_0:jtag_uart_avalon_jtag_slave_address -> jtag_uart:av_address
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_read;                          // mm_interconnect_0:jtag_uart_avalon_jtag_slave_read -> jtag_uart:av_read_n
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_write;                         // mm_interconnect_0:jtag_uart_avalon_jtag_slave_write -> jtag_uart:av_write_n
	wire  [31:0] mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata;                     // mm_interconnect_0:jtag_uart_avalon_jtag_slave_writedata -> jtag_uart:av_writedata
	wire  [31:0] mm_interconnect_0_sysid_qsys_control_slave_readdata;                         // sysid_qsys:readdata -> mm_interconnect_0:sysid_qsys_control_slave_readdata
	wire   [0:0] mm_interconnect_0_sysid_qsys_control_slave_address;                          // mm_interconnect_0:sysid_qsys_control_slave_address -> sysid_qsys:address
	wire  [31:0] mm_interconnect_0_nios2_cpu_debug_mem_slave_readdata;                        // nios2_cpu:debug_mem_slave_readdata -> mm_interconnect_0:nios2_cpu_debug_mem_slave_readdata
	wire         mm_interconnect_0_nios2_cpu_debug_mem_slave_waitrequest;                     // nios2_cpu:debug_mem_slave_waitrequest -> mm_interconnect_0:nios2_cpu_debug_mem_slave_waitrequest
	wire         mm_interconnect_0_nios2_cpu_debug_mem_slave_debugaccess;                     // mm_interconnect_0:nios2_cpu_debug_mem_slave_debugaccess -> nios2_cpu:debug_mem_slave_debugaccess
	wire   [8:0] mm_interconnect_0_nios2_cpu_debug_mem_slave_address;                         // mm_interconnect_0:nios2_cpu_debug_mem_slave_address -> nios2_cpu:debug_mem_slave_address
	wire         mm_interconnect_0_nios2_cpu_debug_mem_slave_read;                            // mm_interconnect_0:nios2_cpu_debug_mem_slave_read -> nios2_cpu:debug_mem_slave_read
	wire   [3:0] mm_interconnect_0_nios2_cpu_debug_mem_slave_byteenable;                      // mm_interconnect_0:nios2_cpu_debug_mem_slave_byteenable -> nios2_cpu:debug_mem_slave_byteenable
	wire         mm_interconnect_0_nios2_cpu_debug_mem_slave_write;                           // mm_interconnect_0:nios2_cpu_debug_mem_slave_write -> nios2_cpu:debug_mem_slave_write
	wire  [31:0] mm_interconnect_0_nios2_cpu_debug_mem_slave_writedata;                       // mm_interconnect_0:nios2_cpu_debug_mem_slave_writedata -> nios2_cpu:debug_mem_slave_writedata
	wire         mm_interconnect_0_onchip_memory2_s1_chipselect;                              // mm_interconnect_0:onchip_memory2_s1_chipselect -> onchip_memory2:chipselect
	wire  [31:0] mm_interconnect_0_onchip_memory2_s1_readdata;                                // onchip_memory2:readdata -> mm_interconnect_0:onchip_memory2_s1_readdata
	wire  [14:0] mm_interconnect_0_onchip_memory2_s1_address;                                 // mm_interconnect_0:onchip_memory2_s1_address -> onchip_memory2:address
	wire   [3:0] mm_interconnect_0_onchip_memory2_s1_byteenable;                              // mm_interconnect_0:onchip_memory2_s1_byteenable -> onchip_memory2:byteenable
	wire         mm_interconnect_0_onchip_memory2_s1_write;                                   // mm_interconnect_0:onchip_memory2_s1_write -> onchip_memory2:write
	wire  [31:0] mm_interconnect_0_onchip_memory2_s1_writedata;                               // mm_interconnect_0:onchip_memory2_s1_writedata -> onchip_memory2:writedata
	wire         mm_interconnect_0_onchip_memory2_s1_clken;                                   // mm_interconnect_0:onchip_memory2_s1_clken -> onchip_memory2:clken
	wire         mm_interconnect_0_sdram_controller_s1_chipselect;                            // mm_interconnect_0:sdram_controller_s1_chipselect -> sdram_controller:az_cs
	wire  [31:0] mm_interconnect_0_sdram_controller_s1_readdata;                              // sdram_controller:za_data -> mm_interconnect_0:sdram_controller_s1_readdata
	wire         mm_interconnect_0_sdram_controller_s1_waitrequest;                           // sdram_controller:za_waitrequest -> mm_interconnect_0:sdram_controller_s1_waitrequest
	wire  [24:0] mm_interconnect_0_sdram_controller_s1_address;                               // mm_interconnect_0:sdram_controller_s1_address -> sdram_controller:az_addr
	wire         mm_interconnect_0_sdram_controller_s1_read;                                  // mm_interconnect_0:sdram_controller_s1_read -> sdram_controller:az_rd_n
	wire   [3:0] mm_interconnect_0_sdram_controller_s1_byteenable;                            // mm_interconnect_0:sdram_controller_s1_byteenable -> sdram_controller:az_be_n
	wire         mm_interconnect_0_sdram_controller_s1_readdatavalid;                         // sdram_controller:za_valid -> mm_interconnect_0:sdram_controller_s1_readdatavalid
	wire         mm_interconnect_0_sdram_controller_s1_write;                                 // mm_interconnect_0:sdram_controller_s1_write -> sdram_controller:az_wr_n
	wire  [31:0] mm_interconnect_0_sdram_controller_s1_writedata;                             // mm_interconnect_0:sdram_controller_s1_writedata -> sdram_controller:az_data
	wire         mm_interconnect_0_pio_touch_s1_chipselect;                                   // mm_interconnect_0:pio_touch_s1_chipselect -> pio_touch:chipselect
	wire  [31:0] mm_interconnect_0_pio_touch_s1_readdata;                                     // pio_touch:readdata -> mm_interconnect_0:pio_touch_s1_readdata
	wire   [1:0] mm_interconnect_0_pio_touch_s1_address;                                      // mm_interconnect_0:pio_touch_s1_address -> pio_touch:address
	wire         mm_interconnect_0_pio_touch_s1_write;                                        // mm_interconnect_0:pio_touch_s1_write -> pio_touch:write_n
	wire  [31:0] mm_interconnect_0_pio_touch_s1_writedata;                                    // mm_interconnect_0:pio_touch_s1_writedata -> pio_touch:writedata
	wire         mm_interconnect_0_timer_s1_chipselect;                                       // mm_interconnect_0:timer_s1_chipselect -> timer:chipselect
	wire  [15:0] mm_interconnect_0_timer_s1_readdata;                                         // timer:readdata -> mm_interconnect_0:timer_s1_readdata
	wire   [2:0] mm_interconnect_0_timer_s1_address;                                          // mm_interconnect_0:timer_s1_address -> timer:address
	wire         mm_interconnect_0_timer_s1_write;                                            // mm_interconnect_0:timer_s1_write -> timer:write_n
	wire  [15:0] mm_interconnect_0_timer_s1_writedata;                                        // mm_interconnect_0:timer_s1_writedata -> timer:writedata
	wire         mm_interconnect_0_spi_touch_spi_control_port_chipselect;                     // mm_interconnect_0:spi_touch_spi_control_port_chipselect -> spi_touch:spi_select
	wire  [15:0] mm_interconnect_0_spi_touch_spi_control_port_readdata;                       // spi_touch:data_to_cpu -> mm_interconnect_0:spi_touch_spi_control_port_readdata
	wire   [2:0] mm_interconnect_0_spi_touch_spi_control_port_address;                        // mm_interconnect_0:spi_touch_spi_control_port_address -> spi_touch:mem_addr
	wire         mm_interconnect_0_spi_touch_spi_control_port_read;                           // mm_interconnect_0:spi_touch_spi_control_port_read -> spi_touch:read_n
	wire         mm_interconnect_0_spi_touch_spi_control_port_write;                          // mm_interconnect_0:spi_touch_spi_control_port_write -> spi_touch:write_n
	wire  [15:0] mm_interconnect_0_spi_touch_spi_control_port_writedata;                      // mm_interconnect_0:spi_touch_spi_control_port_writedata -> spi_touch:data_from_cpu
	wire         irq_mapper_receiver1_irq;                                                    // jtag_uart:av_irq -> irq_mapper:receiver1_irq
	wire         irq_mapper_receiver2_irq;                                                    // pio_touch:irq -> irq_mapper:receiver2_irq
	wire         irq_mapper_receiver3_irq;                                                    // timer:irq -> irq_mapper:receiver3_irq
	wire  [31:0] nios2_cpu_irq_irq;                                                           // irq_mapper:sender_irq -> nios2_cpu:irq
	wire         irq_mapper_receiver0_irq;                                                    // irq_synchronizer:sender_irq -> irq_mapper:receiver0_irq
	wire   [0:0] irq_synchronizer_receiver_irq;                                               // audio:irq -> irq_synchronizer:receiver_irq
	wire         rst_controller_reset_out_reset;                                              // rst_controller:reset_out -> [audio:reset, audio_and_video_config:reset, irq_synchronizer:receiver_reset, mm_interconnect_0:audio_reset_reset_bridge_in_reset_reset]
	wire         nios2_cpu_debug_reset_request_reset;                                         // nios2_cpu:debug_reset_request -> [rst_controller:reset_in1, rst_controller_002:reset_in1, rst_controller_004:reset_in1, rst_controller_005:reset_in0]
	wire         audio_pll_reset_source_reset;                                                // audio_pll:reset_source_reset -> rst_controller:reset_in2
	wire         rst_controller_001_reset_out_reset;                                          // rst_controller_001:reset_out -> [audio_pll:ref_reset_reset, video_pll:ref_reset_reset]
	wire         rst_controller_002_reset_out_reset;                                          // rst_controller_002:reset_out -> [irq_mapper:reset, irq_synchronizer:sender_reset, jtag_uart:rst_n, mm_interconnect_0:video_pixel_buffer_dma_reset_reset_bridge_in_reset_reset, nios2_cpu:reset_n, onchip_memory2:reset, pio_touch:reset_n, rst_translator:in_reset, sdram_controller:reset_n, spi_touch:reset_n, sram:reset, sysid_qsys:reset_n, video_pixel_buffer_dma:reset, video_rgb_resampler_0:reset]
	wire         rst_controller_002_reset_out_reset_req;                                      // rst_controller_002:reset_req -> [nios2_cpu:reset_req, onchip_memory2:reset_req, rst_translator:reset_req_in]
	wire         sys_sdram_pll_reset_source_reset;                                            // sys_sdram_pll:reset_source_reset -> [rst_controller_002:reset_in2, rst_controller_005:reset_in1]
	wire         rst_controller_003_reset_out_reset;                                          // rst_controller_003:reset_out -> sys_sdram_pll:ref_reset_reset
	wire         rst_controller_004_reset_out_reset;                                          // rst_controller_004:reset_out -> [mm_interconnect_0:timer_reset_reset_bridge_in_reset_reset, timer:reset_n]
	wire         rst_controller_005_reset_out_reset;                                          // rst_controller_005:reset_out -> video_dual_clock_buffer:reset_stream_in
	wire         rst_controller_006_reset_out_reset;                                          // rst_controller_006:reset_out -> video_dual_clock_buffer:reset_stream_out
	wire         video_pll_reset_source_reset;                                                // video_pll:reset_source_reset -> [rst_controller_006:reset_in0, rst_controller_007:reset_in1]
	wire         rst_controller_007_reset_out_reset;                                          // rst_controller_007:reset_out -> video_vga_controller:reset

	Core_audio audio (
		.clk         (clock_bridge_out_clk_clk),                              //                clk.clk
		.reset       (rst_controller_reset_out_reset),                        //              reset.reset
		.address     (mm_interconnect_0_audio_avalon_audio_slave_address),    // avalon_audio_slave.address
		.chipselect  (mm_interconnect_0_audio_avalon_audio_slave_chipselect), //                   .chipselect
		.read        (mm_interconnect_0_audio_avalon_audio_slave_read),       //                   .read
		.write       (mm_interconnect_0_audio_avalon_audio_slave_write),      //                   .write
		.writedata   (mm_interconnect_0_audio_avalon_audio_slave_writedata),  //                   .writedata
		.readdata    (mm_interconnect_0_audio_avalon_audio_slave_readdata),   //                   .readdata
		.irq         (irq_synchronizer_receiver_irq),                         //          interrupt.irq
		.AUD_ADCDAT  (audio_external_interface_ADCDAT),                       // external_interface.export
		.AUD_ADCLRCK (audio_external_interface_ADCLRCK),                      //                   .export
		.AUD_BCLK    (audio_external_interface_BCLK),                         //                   .export
		.AUD_DACDAT  (audio_external_interface_DACDAT),                       //                   .export
		.AUD_DACLRCK (audio_external_interface_DACLRCK)                       //                   .export
	);

	Core_audio_and_video_config audio_and_video_config (
		.clk         (clock_bridge_out_clk_clk),                                                    //                    clk.clk
		.reset       (rst_controller_reset_out_reset),                                              //                  reset.reset
		.address     (mm_interconnect_0_audio_and_video_config_avalon_av_config_slave_address),     // avalon_av_config_slave.address
		.byteenable  (mm_interconnect_0_audio_and_video_config_avalon_av_config_slave_byteenable),  //                       .byteenable
		.read        (mm_interconnect_0_audio_and_video_config_avalon_av_config_slave_read),        //                       .read
		.write       (mm_interconnect_0_audio_and_video_config_avalon_av_config_slave_write),       //                       .write
		.writedata   (mm_interconnect_0_audio_and_video_config_avalon_av_config_slave_writedata),   //                       .writedata
		.readdata    (mm_interconnect_0_audio_and_video_config_avalon_av_config_slave_readdata),    //                       .readdata
		.waitrequest (mm_interconnect_0_audio_and_video_config_avalon_av_config_slave_waitrequest), //                       .waitrequest
		.I2C_SDAT    (audio_and_video_config_external_interface_SDAT),                              //     external_interface.export
		.I2C_SCLK    (audio_and_video_config_external_interface_SCLK)                               //                       .export
	);

	Core_audio_pll audio_pll (
		.ref_clk_clk        (clk_clk),                            //      ref_clk.clk
		.ref_reset_reset    (rst_controller_001_reset_out_reset), //    ref_reset.reset
		.audio_clk_clk      (clock_bridge_out_clk_clk),           //    audio_clk.clk
		.reset_source_reset (audio_pll_reset_source_reset)        // reset_source.reset
	);

	Core_jtag_uart jtag_uart (
		.clk            (sys_sdram_pll_sys_clk_clk),                                 //               clk.clk
		.rst_n          (~rst_controller_002_reset_out_reset),                       //             reset.reset_n
		.av_chipselect  (mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (mm_interconnect_0_jtag_uart_avalon_jtag_slave_address),     //                  .address
		.av_read_n      (~mm_interconnect_0_jtag_uart_avalon_jtag_slave_read),       //                  .read_n
		.av_readdata    (mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata),    //                  .readdata
		.av_write_n     (~mm_interconnect_0_jtag_uart_avalon_jtag_slave_write),      //                  .write_n
		.av_writedata   (mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata),   //                  .writedata
		.av_waitrequest (mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest), //                  .waitrequest
		.av_irq         (irq_mapper_receiver1_irq)                                   //               irq.irq
	);

	Core_nios2_cpu nios2_cpu (
		.clk                                 (sys_sdram_pll_sys_clk_clk),                               //                       clk.clk
		.reset_n                             (~rst_controller_002_reset_out_reset),                     //                     reset.reset_n
		.reset_req                           (rst_controller_002_reset_out_reset_req),                  //                          .reset_req
		.d_address                           (nios2_cpu_data_master_address),                           //               data_master.address
		.d_byteenable                        (nios2_cpu_data_master_byteenable),                        //                          .byteenable
		.d_read                              (nios2_cpu_data_master_read),                              //                          .read
		.d_readdata                          (nios2_cpu_data_master_readdata),                          //                          .readdata
		.d_waitrequest                       (nios2_cpu_data_master_waitrequest),                       //                          .waitrequest
		.d_write                             (nios2_cpu_data_master_write),                             //                          .write
		.d_writedata                         (nios2_cpu_data_master_writedata),                         //                          .writedata
		.d_readdatavalid                     (nios2_cpu_data_master_readdatavalid),                     //                          .readdatavalid
		.debug_mem_slave_debugaccess_to_roms (nios2_cpu_data_master_debugaccess),                       //                          .debugaccess
		.i_address                           (nios2_cpu_instruction_master_address),                    //        instruction_master.address
		.i_read                              (nios2_cpu_instruction_master_read),                       //                          .read
		.i_readdata                          (nios2_cpu_instruction_master_readdata),                   //                          .readdata
		.i_waitrequest                       (nios2_cpu_instruction_master_waitrequest),                //                          .waitrequest
		.i_readdatavalid                     (nios2_cpu_instruction_master_readdatavalid),              //                          .readdatavalid
		.irq                                 (nios2_cpu_irq_irq),                                       //                       irq.irq
		.debug_reset_request                 (nios2_cpu_debug_reset_request_reset),                     //       debug_reset_request.reset
		.debug_mem_slave_address             (mm_interconnect_0_nios2_cpu_debug_mem_slave_address),     //           debug_mem_slave.address
		.debug_mem_slave_byteenable          (mm_interconnect_0_nios2_cpu_debug_mem_slave_byteenable),  //                          .byteenable
		.debug_mem_slave_debugaccess         (mm_interconnect_0_nios2_cpu_debug_mem_slave_debugaccess), //                          .debugaccess
		.debug_mem_slave_read                (mm_interconnect_0_nios2_cpu_debug_mem_slave_read),        //                          .read
		.debug_mem_slave_readdata            (mm_interconnect_0_nios2_cpu_debug_mem_slave_readdata),    //                          .readdata
		.debug_mem_slave_waitrequest         (mm_interconnect_0_nios2_cpu_debug_mem_slave_waitrequest), //                          .waitrequest
		.debug_mem_slave_write               (mm_interconnect_0_nios2_cpu_debug_mem_slave_write),       //                          .write
		.debug_mem_slave_writedata           (mm_interconnect_0_nios2_cpu_debug_mem_slave_writedata),   //                          .writedata
		.dummy_ci_port                       ()                                                         // custom_instruction_master.readra
	);

	Core_onchip_memory2 onchip_memory2 (
		.clk        (sys_sdram_pll_sys_clk_clk),                      //   clk1.clk
		.address    (mm_interconnect_0_onchip_memory2_s1_address),    //     s1.address
		.clken      (mm_interconnect_0_onchip_memory2_s1_clken),      //       .clken
		.chipselect (mm_interconnect_0_onchip_memory2_s1_chipselect), //       .chipselect
		.write      (mm_interconnect_0_onchip_memory2_s1_write),      //       .write
		.readdata   (mm_interconnect_0_onchip_memory2_s1_readdata),   //       .readdata
		.writedata  (mm_interconnect_0_onchip_memory2_s1_writedata),  //       .writedata
		.byteenable (mm_interconnect_0_onchip_memory2_s1_byteenable), //       .byteenable
		.reset      (rst_controller_002_reset_out_reset),             // reset1.reset
		.reset_req  (rst_controller_002_reset_out_reset_req)          //       .reset_req
	);

	Core_pio_touch pio_touch (
		.clk        (sys_sdram_pll_sys_clk_clk),                 //                 clk.clk
		.reset_n    (~rst_controller_002_reset_out_reset),       //               reset.reset_n
		.address    (mm_interconnect_0_pio_touch_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_pio_touch_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_pio_touch_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_pio_touch_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_pio_touch_s1_readdata),   //                    .readdata
		.in_port    (pio_touch_external_connection_export),      // external_connection.export
		.irq        (irq_mapper_receiver2_irq)                   //                 irq.irq
	);

	Core_sdram_controller sdram_controller (
		.clk            (sys_sdram_pll_sys_clk_clk),                           //   clk.clk
		.reset_n        (~rst_controller_002_reset_out_reset),                 // reset.reset_n
		.az_addr        (mm_interconnect_0_sdram_controller_s1_address),       //    s1.address
		.az_be_n        (~mm_interconnect_0_sdram_controller_s1_byteenable),   //      .byteenable_n
		.az_cs          (mm_interconnect_0_sdram_controller_s1_chipselect),    //      .chipselect
		.az_data        (mm_interconnect_0_sdram_controller_s1_writedata),     //      .writedata
		.az_rd_n        (~mm_interconnect_0_sdram_controller_s1_read),         //      .read_n
		.az_wr_n        (~mm_interconnect_0_sdram_controller_s1_write),        //      .write_n
		.za_data        (mm_interconnect_0_sdram_controller_s1_readdata),      //      .readdata
		.za_valid       (mm_interconnect_0_sdram_controller_s1_readdatavalid), //      .readdatavalid
		.za_waitrequest (mm_interconnect_0_sdram_controller_s1_waitrequest),   //      .waitrequest
		.zs_addr        (sdram_controller_wire_addr),                          //  wire.export
		.zs_ba          (sdram_controller_wire_ba),                            //      .export
		.zs_cas_n       (sdram_controller_wire_cas_n),                         //      .export
		.zs_cke         (sdram_controller_wire_cke),                           //      .export
		.zs_cs_n        (sdram_controller_wire_cs_n),                          //      .export
		.zs_dq          (sdram_controller_wire_dq),                            //      .export
		.zs_dqm         (sdram_controller_wire_dqm),                           //      .export
		.zs_ras_n       (sdram_controller_wire_ras_n),                         //      .export
		.zs_we_n        (sdram_controller_wire_we_n)                           //      .export
	);

	Core_spi_touch spi_touch (
		.clk           (sys_sdram_pll_sys_clk_clk),                               //              clk.clk
		.reset_n       (~rst_controller_002_reset_out_reset),                     //            reset.reset_n
		.data_from_cpu (mm_interconnect_0_spi_touch_spi_control_port_writedata),  // spi_control_port.writedata
		.data_to_cpu   (mm_interconnect_0_spi_touch_spi_control_port_readdata),   //                 .readdata
		.mem_addr      (mm_interconnect_0_spi_touch_spi_control_port_address),    //                 .address
		.read_n        (~mm_interconnect_0_spi_touch_spi_control_port_read),      //                 .read_n
		.spi_select    (mm_interconnect_0_spi_touch_spi_control_port_chipselect), //                 .chipselect
		.write_n       (~mm_interconnect_0_spi_touch_spi_control_port_write),     //                 .write_n
		.irq           (),                                                        //              irq.irq
		.MISO          (spi_touch_external_MISO),                                 //         external.export
		.MOSI          (spi_touch_external_MOSI),                                 //                 .export
		.SCLK          (spi_touch_external_SCLK),                                 //                 .export
		.SS_n          (spi_touch_external_SS_n)                                  //                 .export
	);

	Core_sram sram (
		.clk           (sys_sdram_pll_sys_clk_clk),                              //                clk.clk
		.reset         (rst_controller_002_reset_out_reset),                     //              reset.reset
		.SRAM_DQ       (sram_external_interface_DQ),                             // external_interface.export
		.SRAM_ADDR     (sram_external_interface_ADDR),                           //                   .export
		.SRAM_LB_N     (sram_external_interface_LB_N),                           //                   .export
		.SRAM_UB_N     (sram_external_interface_UB_N),                           //                   .export
		.SRAM_CE_N     (sram_external_interface_CE_N),                           //                   .export
		.SRAM_OE_N     (sram_external_interface_OE_N),                           //                   .export
		.SRAM_WE_N     (sram_external_interface_WE_N),                           //                   .export
		.address       (mm_interconnect_0_sram_avalon_sram_slave_address),       //  avalon_sram_slave.address
		.byteenable    (mm_interconnect_0_sram_avalon_sram_slave_byteenable),    //                   .byteenable
		.read          (mm_interconnect_0_sram_avalon_sram_slave_read),          //                   .read
		.write         (mm_interconnect_0_sram_avalon_sram_slave_write),         //                   .write
		.writedata     (mm_interconnect_0_sram_avalon_sram_slave_writedata),     //                   .writedata
		.readdata      (mm_interconnect_0_sram_avalon_sram_slave_readdata),      //                   .readdata
		.readdatavalid (mm_interconnect_0_sram_avalon_sram_slave_readdatavalid)  //                   .readdatavalid
	);

	Core_sys_sdram_pll sys_sdram_pll (
		.ref_clk_clk        (clk_0_clk),                          //      ref_clk.clk
		.ref_reset_reset    (rst_controller_003_reset_out_reset), //    ref_reset.reset
		.sys_clk_clk        (sys_sdram_pll_sys_clk_clk),          //      sys_clk.clk
		.sdram_clk_clk      (sys_sdram_pll_sdram_clk_clk),        //    sdram_clk.clk
		.reset_source_reset (sys_sdram_pll_reset_source_reset)    // reset_source.reset
	);

	Core_sysid_qsys sysid_qsys (
		.clock    (sys_sdram_pll_sys_clk_clk),                           //           clk.clk
		.reset_n  (~rst_controller_002_reset_out_reset),                 //         reset.reset_n
		.readdata (mm_interconnect_0_sysid_qsys_control_slave_readdata), // control_slave.readdata
		.address  (mm_interconnect_0_sysid_qsys_control_slave_address)   //              .address
	);

	Core_timer timer (
		.clk        (sys_sdram_pll_sys_clk_clk),             //   clk.clk
		.reset_n    (~rst_controller_004_reset_out_reset),   // reset.reset_n
		.address    (mm_interconnect_0_timer_s1_address),    //    s1.address
		.writedata  (mm_interconnect_0_timer_s1_writedata),  //      .writedata
		.readdata   (mm_interconnect_0_timer_s1_readdata),   //      .readdata
		.chipselect (mm_interconnect_0_timer_s1_chipselect), //      .chipselect
		.write_n    (~mm_interconnect_0_timer_s1_write),     //      .write_n
		.irq        (irq_mapper_receiver3_irq)               //   irq.irq
	);

	Core_video_dual_clock_buffer video_dual_clock_buffer (
		.clk_stream_in            (sys_sdram_pll_sys_clk_clk),                                     //         clock_stream_in.clk
		.reset_stream_in          (rst_controller_005_reset_out_reset),                            //         reset_stream_in.reset
		.clk_stream_out           (video_pll_lcd_clk_clk),                                         //        clock_stream_out.clk
		.reset_stream_out         (rst_controller_006_reset_out_reset),                            //        reset_stream_out.reset
		.stream_in_ready          (video_rgb_resampler_0_avalon_rgb_source_ready),                 //   avalon_dc_buffer_sink.ready
		.stream_in_startofpacket  (video_rgb_resampler_0_avalon_rgb_source_startofpacket),         //                        .startofpacket
		.stream_in_endofpacket    (video_rgb_resampler_0_avalon_rgb_source_endofpacket),           //                        .endofpacket
		.stream_in_valid          (video_rgb_resampler_0_avalon_rgb_source_valid),                 //                        .valid
		.stream_in_data           (video_rgb_resampler_0_avalon_rgb_source_data),                  //                        .data
		.stream_out_ready         (video_dual_clock_buffer_avalon_dc_buffer_source_ready),         // avalon_dc_buffer_source.ready
		.stream_out_startofpacket (video_dual_clock_buffer_avalon_dc_buffer_source_startofpacket), //                        .startofpacket
		.stream_out_endofpacket   (video_dual_clock_buffer_avalon_dc_buffer_source_endofpacket),   //                        .endofpacket
		.stream_out_valid         (video_dual_clock_buffer_avalon_dc_buffer_source_valid),         //                        .valid
		.stream_out_data          (video_dual_clock_buffer_avalon_dc_buffer_source_data)           //                        .data
	);

	Core_video_pixel_buffer_dma video_pixel_buffer_dma (
		.clk                  (sys_sdram_pll_sys_clk_clk),                                                //                     clk.clk
		.reset                (rst_controller_002_reset_out_reset),                                       //                   reset.reset
		.master_readdatavalid (video_pixel_buffer_dma_avalon_pixel_dma_master_readdatavalid),             // avalon_pixel_dma_master.readdatavalid
		.master_waitrequest   (video_pixel_buffer_dma_avalon_pixel_dma_master_waitrequest),               //                        .waitrequest
		.master_address       (video_pixel_buffer_dma_avalon_pixel_dma_master_address),                   //                        .address
		.master_arbiterlock   (video_pixel_buffer_dma_avalon_pixel_dma_master_lock),                      //                        .lock
		.master_read          (video_pixel_buffer_dma_avalon_pixel_dma_master_read),                      //                        .read
		.master_readdata      (video_pixel_buffer_dma_avalon_pixel_dma_master_readdata),                  //                        .readdata
		.slave_address        (mm_interconnect_0_video_pixel_buffer_dma_avalon_control_slave_address),    //    avalon_control_slave.address
		.slave_byteenable     (mm_interconnect_0_video_pixel_buffer_dma_avalon_control_slave_byteenable), //                        .byteenable
		.slave_read           (mm_interconnect_0_video_pixel_buffer_dma_avalon_control_slave_read),       //                        .read
		.slave_write          (mm_interconnect_0_video_pixel_buffer_dma_avalon_control_slave_write),      //                        .write
		.slave_writedata      (mm_interconnect_0_video_pixel_buffer_dma_avalon_control_slave_writedata),  //                        .writedata
		.slave_readdata       (mm_interconnect_0_video_pixel_buffer_dma_avalon_control_slave_readdata),   //                        .readdata
		.stream_ready         (video_pixel_buffer_dma_avalon_pixel_source_ready),                         //     avalon_pixel_source.ready
		.stream_startofpacket (video_pixel_buffer_dma_avalon_pixel_source_startofpacket),                 //                        .startofpacket
		.stream_endofpacket   (video_pixel_buffer_dma_avalon_pixel_source_endofpacket),                   //                        .endofpacket
		.stream_valid         (video_pixel_buffer_dma_avalon_pixel_source_valid),                         //                        .valid
		.stream_data          (video_pixel_buffer_dma_avalon_pixel_source_data)                           //                        .data
	);

	Core_video_pll video_pll (
		.ref_clk_clk        (clk_clk),                            //      ref_clk.clk
		.ref_reset_reset    (rst_controller_001_reset_out_reset), //    ref_reset.reset
		.lcd_clk_clk        (video_pll_lcd_clk_clk),              //      lcd_clk.clk
		.reset_source_reset (video_pll_reset_source_reset)        // reset_source.reset
	);

	Core_video_rgb_resampler_0 video_rgb_resampler_0 (
		.clk                      (sys_sdram_pll_sys_clk_clk),                                //               clk.clk
		.reset                    (rst_controller_002_reset_out_reset),                       //             reset.reset
		.stream_in_startofpacket  (video_pixel_buffer_dma_avalon_pixel_source_startofpacket), //   avalon_rgb_sink.startofpacket
		.stream_in_endofpacket    (video_pixel_buffer_dma_avalon_pixel_source_endofpacket),   //                  .endofpacket
		.stream_in_valid          (video_pixel_buffer_dma_avalon_pixel_source_valid),         //                  .valid
		.stream_in_ready          (video_pixel_buffer_dma_avalon_pixel_source_ready),         //                  .ready
		.stream_in_data           (video_pixel_buffer_dma_avalon_pixel_source_data),          //                  .data
		.stream_out_ready         (video_rgb_resampler_0_avalon_rgb_source_ready),            // avalon_rgb_source.ready
		.stream_out_startofpacket (video_rgb_resampler_0_avalon_rgb_source_startofpacket),    //                  .startofpacket
		.stream_out_endofpacket   (video_rgb_resampler_0_avalon_rgb_source_endofpacket),      //                  .endofpacket
		.stream_out_valid         (video_rgb_resampler_0_avalon_rgb_source_valid),            //                  .valid
		.stream_out_data          (video_rgb_resampler_0_avalon_rgb_source_data)              //                  .data
	);

	Core_video_vga_controller video_vga_controller (
		.clk           (video_pll_lcd_clk_clk),                                         //                clk.clk
		.reset         (rst_controller_007_reset_out_reset),                            //              reset.reset
		.data          (video_dual_clock_buffer_avalon_dc_buffer_source_data),          //    avalon_vga_sink.data
		.startofpacket (video_dual_clock_buffer_avalon_dc_buffer_source_startofpacket), //                   .startofpacket
		.endofpacket   (video_dual_clock_buffer_avalon_dc_buffer_source_endofpacket),   //                   .endofpacket
		.valid         (video_dual_clock_buffer_avalon_dc_buffer_source_valid),         //                   .valid
		.ready         (video_dual_clock_buffer_avalon_dc_buffer_source_ready),         //                   .ready
		.VGA_CLK       (video_vga_controller_external_interface_CLK),                   // external_interface.export
		.VGA_HS        (video_vga_controller_external_interface_HS),                    //                   .export
		.VGA_VS        (video_vga_controller_external_interface_VS),                    //                   .export
		.VGA_BLANK     (video_vga_controller_external_interface_BLANK),                 //                   .export
		.VGA_SYNC      (video_vga_controller_external_interface_SYNC),                  //                   .export
		.VGA_DATA_EN   (video_vga_controller_external_interface_DATA_EN),               //                   .export
		.VGA_R         (video_vga_controller_external_interface_R),                     //                   .export
		.VGA_G         (video_vga_controller_external_interface_G),                     //                   .export
		.VGA_B         (video_vga_controller_external_interface_B)                      //                   .export
	);

	Core_mm_interconnect_0 mm_interconnect_0 (
		.audio_pll_audio_clk_clk                                      (clock_bridge_out_clk_clk),                                                    //                                audio_pll_audio_clk.clk
		.sys_sdram_pll_sys_clk_clk                                    (sys_sdram_pll_sys_clk_clk),                                                   //                              sys_sdram_pll_sys_clk.clk
		.audio_reset_reset_bridge_in_reset_reset                      (rst_controller_reset_out_reset),                                              //                  audio_reset_reset_bridge_in_reset.reset
		.timer_reset_reset_bridge_in_reset_reset                      (rst_controller_004_reset_out_reset),                                          //                  timer_reset_reset_bridge_in_reset.reset
		.video_pixel_buffer_dma_reset_reset_bridge_in_reset_reset     (rst_controller_002_reset_out_reset),                                          // video_pixel_buffer_dma_reset_reset_bridge_in_reset.reset
		.nios2_cpu_data_master_address                                (nios2_cpu_data_master_address),                                               //                              nios2_cpu_data_master.address
		.nios2_cpu_data_master_waitrequest                            (nios2_cpu_data_master_waitrequest),                                           //                                                   .waitrequest
		.nios2_cpu_data_master_byteenable                             (nios2_cpu_data_master_byteenable),                                            //                                                   .byteenable
		.nios2_cpu_data_master_read                                   (nios2_cpu_data_master_read),                                                  //                                                   .read
		.nios2_cpu_data_master_readdata                               (nios2_cpu_data_master_readdata),                                              //                                                   .readdata
		.nios2_cpu_data_master_readdatavalid                          (nios2_cpu_data_master_readdatavalid),                                         //                                                   .readdatavalid
		.nios2_cpu_data_master_write                                  (nios2_cpu_data_master_write),                                                 //                                                   .write
		.nios2_cpu_data_master_writedata                              (nios2_cpu_data_master_writedata),                                             //                                                   .writedata
		.nios2_cpu_data_master_debugaccess                            (nios2_cpu_data_master_debugaccess),                                           //                                                   .debugaccess
		.nios2_cpu_instruction_master_address                         (nios2_cpu_instruction_master_address),                                        //                       nios2_cpu_instruction_master.address
		.nios2_cpu_instruction_master_waitrequest                     (nios2_cpu_instruction_master_waitrequest),                                    //                                                   .waitrequest
		.nios2_cpu_instruction_master_read                            (nios2_cpu_instruction_master_read),                                           //                                                   .read
		.nios2_cpu_instruction_master_readdata                        (nios2_cpu_instruction_master_readdata),                                       //                                                   .readdata
		.nios2_cpu_instruction_master_readdatavalid                   (nios2_cpu_instruction_master_readdatavalid),                                  //                                                   .readdatavalid
		.video_pixel_buffer_dma_avalon_pixel_dma_master_address       (video_pixel_buffer_dma_avalon_pixel_dma_master_address),                      //     video_pixel_buffer_dma_avalon_pixel_dma_master.address
		.video_pixel_buffer_dma_avalon_pixel_dma_master_waitrequest   (video_pixel_buffer_dma_avalon_pixel_dma_master_waitrequest),                  //                                                   .waitrequest
		.video_pixel_buffer_dma_avalon_pixel_dma_master_read          (video_pixel_buffer_dma_avalon_pixel_dma_master_read),                         //                                                   .read
		.video_pixel_buffer_dma_avalon_pixel_dma_master_readdata      (video_pixel_buffer_dma_avalon_pixel_dma_master_readdata),                     //                                                   .readdata
		.video_pixel_buffer_dma_avalon_pixel_dma_master_readdatavalid (video_pixel_buffer_dma_avalon_pixel_dma_master_readdatavalid),                //                                                   .readdatavalid
		.video_pixel_buffer_dma_avalon_pixel_dma_master_lock          (video_pixel_buffer_dma_avalon_pixel_dma_master_lock),                         //                                                   .lock
		.audio_avalon_audio_slave_address                             (mm_interconnect_0_audio_avalon_audio_slave_address),                          //                           audio_avalon_audio_slave.address
		.audio_avalon_audio_slave_write                               (mm_interconnect_0_audio_avalon_audio_slave_write),                            //                                                   .write
		.audio_avalon_audio_slave_read                                (mm_interconnect_0_audio_avalon_audio_slave_read),                             //                                                   .read
		.audio_avalon_audio_slave_readdata                            (mm_interconnect_0_audio_avalon_audio_slave_readdata),                         //                                                   .readdata
		.audio_avalon_audio_slave_writedata                           (mm_interconnect_0_audio_avalon_audio_slave_writedata),                        //                                                   .writedata
		.audio_avalon_audio_slave_chipselect                          (mm_interconnect_0_audio_avalon_audio_slave_chipselect),                       //                                                   .chipselect
		.audio_and_video_config_avalon_av_config_slave_address        (mm_interconnect_0_audio_and_video_config_avalon_av_config_slave_address),     //      audio_and_video_config_avalon_av_config_slave.address
		.audio_and_video_config_avalon_av_config_slave_write          (mm_interconnect_0_audio_and_video_config_avalon_av_config_slave_write),       //                                                   .write
		.audio_and_video_config_avalon_av_config_slave_read           (mm_interconnect_0_audio_and_video_config_avalon_av_config_slave_read),        //                                                   .read
		.audio_and_video_config_avalon_av_config_slave_readdata       (mm_interconnect_0_audio_and_video_config_avalon_av_config_slave_readdata),    //                                                   .readdata
		.audio_and_video_config_avalon_av_config_slave_writedata      (mm_interconnect_0_audio_and_video_config_avalon_av_config_slave_writedata),   //                                                   .writedata
		.audio_and_video_config_avalon_av_config_slave_byteenable     (mm_interconnect_0_audio_and_video_config_avalon_av_config_slave_byteenable),  //                                                   .byteenable
		.audio_and_video_config_avalon_av_config_slave_waitrequest    (mm_interconnect_0_audio_and_video_config_avalon_av_config_slave_waitrequest), //                                                   .waitrequest
		.jtag_uart_avalon_jtag_slave_address                          (mm_interconnect_0_jtag_uart_avalon_jtag_slave_address),                       //                        jtag_uart_avalon_jtag_slave.address
		.jtag_uart_avalon_jtag_slave_write                            (mm_interconnect_0_jtag_uart_avalon_jtag_slave_write),                         //                                                   .write
		.jtag_uart_avalon_jtag_slave_read                             (mm_interconnect_0_jtag_uart_avalon_jtag_slave_read),                          //                                                   .read
		.jtag_uart_avalon_jtag_slave_readdata                         (mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata),                      //                                                   .readdata
		.jtag_uart_avalon_jtag_slave_writedata                        (mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata),                     //                                                   .writedata
		.jtag_uart_avalon_jtag_slave_waitrequest                      (mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest),                   //                                                   .waitrequest
		.jtag_uart_avalon_jtag_slave_chipselect                       (mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect),                    //                                                   .chipselect
		.nios2_cpu_debug_mem_slave_address                            (mm_interconnect_0_nios2_cpu_debug_mem_slave_address),                         //                          nios2_cpu_debug_mem_slave.address
		.nios2_cpu_debug_mem_slave_write                              (mm_interconnect_0_nios2_cpu_debug_mem_slave_write),                           //                                                   .write
		.nios2_cpu_debug_mem_slave_read                               (mm_interconnect_0_nios2_cpu_debug_mem_slave_read),                            //                                                   .read
		.nios2_cpu_debug_mem_slave_readdata                           (mm_interconnect_0_nios2_cpu_debug_mem_slave_readdata),                        //                                                   .readdata
		.nios2_cpu_debug_mem_slave_writedata                          (mm_interconnect_0_nios2_cpu_debug_mem_slave_writedata),                       //                                                   .writedata
		.nios2_cpu_debug_mem_slave_byteenable                         (mm_interconnect_0_nios2_cpu_debug_mem_slave_byteenable),                      //                                                   .byteenable
		.nios2_cpu_debug_mem_slave_waitrequest                        (mm_interconnect_0_nios2_cpu_debug_mem_slave_waitrequest),                     //                                                   .waitrequest
		.nios2_cpu_debug_mem_slave_debugaccess                        (mm_interconnect_0_nios2_cpu_debug_mem_slave_debugaccess),                     //                                                   .debugaccess
		.onchip_memory2_s1_address                                    (mm_interconnect_0_onchip_memory2_s1_address),                                 //                                  onchip_memory2_s1.address
		.onchip_memory2_s1_write                                      (mm_interconnect_0_onchip_memory2_s1_write),                                   //                                                   .write
		.onchip_memory2_s1_readdata                                   (mm_interconnect_0_onchip_memory2_s1_readdata),                                //                                                   .readdata
		.onchip_memory2_s1_writedata                                  (mm_interconnect_0_onchip_memory2_s1_writedata),                               //                                                   .writedata
		.onchip_memory2_s1_byteenable                                 (mm_interconnect_0_onchip_memory2_s1_byteenable),                              //                                                   .byteenable
		.onchip_memory2_s1_chipselect                                 (mm_interconnect_0_onchip_memory2_s1_chipselect),                              //                                                   .chipselect
		.onchip_memory2_s1_clken                                      (mm_interconnect_0_onchip_memory2_s1_clken),                                   //                                                   .clken
		.pio_touch_s1_address                                         (mm_interconnect_0_pio_touch_s1_address),                                      //                                       pio_touch_s1.address
		.pio_touch_s1_write                                           (mm_interconnect_0_pio_touch_s1_write),                                        //                                                   .write
		.pio_touch_s1_readdata                                        (mm_interconnect_0_pio_touch_s1_readdata),                                     //                                                   .readdata
		.pio_touch_s1_writedata                                       (mm_interconnect_0_pio_touch_s1_writedata),                                    //                                                   .writedata
		.pio_touch_s1_chipselect                                      (mm_interconnect_0_pio_touch_s1_chipselect),                                   //                                                   .chipselect
		.sdram_controller_s1_address                                  (mm_interconnect_0_sdram_controller_s1_address),                               //                                sdram_controller_s1.address
		.sdram_controller_s1_write                                    (mm_interconnect_0_sdram_controller_s1_write),                                 //                                                   .write
		.sdram_controller_s1_read                                     (mm_interconnect_0_sdram_controller_s1_read),                                  //                                                   .read
		.sdram_controller_s1_readdata                                 (mm_interconnect_0_sdram_controller_s1_readdata),                              //                                                   .readdata
		.sdram_controller_s1_writedata                                (mm_interconnect_0_sdram_controller_s1_writedata),                             //                                                   .writedata
		.sdram_controller_s1_byteenable                               (mm_interconnect_0_sdram_controller_s1_byteenable),                            //                                                   .byteenable
		.sdram_controller_s1_readdatavalid                            (mm_interconnect_0_sdram_controller_s1_readdatavalid),                         //                                                   .readdatavalid
		.sdram_controller_s1_waitrequest                              (mm_interconnect_0_sdram_controller_s1_waitrequest),                           //                                                   .waitrequest
		.sdram_controller_s1_chipselect                               (mm_interconnect_0_sdram_controller_s1_chipselect),                            //                                                   .chipselect
		.spi_touch_spi_control_port_address                           (mm_interconnect_0_spi_touch_spi_control_port_address),                        //                         spi_touch_spi_control_port.address
		.spi_touch_spi_control_port_write                             (mm_interconnect_0_spi_touch_spi_control_port_write),                          //                                                   .write
		.spi_touch_spi_control_port_read                              (mm_interconnect_0_spi_touch_spi_control_port_read),                           //                                                   .read
		.spi_touch_spi_control_port_readdata                          (mm_interconnect_0_spi_touch_spi_control_port_readdata),                       //                                                   .readdata
		.spi_touch_spi_control_port_writedata                         (mm_interconnect_0_spi_touch_spi_control_port_writedata),                      //                                                   .writedata
		.spi_touch_spi_control_port_chipselect                        (mm_interconnect_0_spi_touch_spi_control_port_chipselect),                     //                                                   .chipselect
		.sram_avalon_sram_slave_address                               (mm_interconnect_0_sram_avalon_sram_slave_address),                            //                             sram_avalon_sram_slave.address
		.sram_avalon_sram_slave_write                                 (mm_interconnect_0_sram_avalon_sram_slave_write),                              //                                                   .write
		.sram_avalon_sram_slave_read                                  (mm_interconnect_0_sram_avalon_sram_slave_read),                               //                                                   .read
		.sram_avalon_sram_slave_readdata                              (mm_interconnect_0_sram_avalon_sram_slave_readdata),                           //                                                   .readdata
		.sram_avalon_sram_slave_writedata                             (mm_interconnect_0_sram_avalon_sram_slave_writedata),                          //                                                   .writedata
		.sram_avalon_sram_slave_byteenable                            (mm_interconnect_0_sram_avalon_sram_slave_byteenable),                         //                                                   .byteenable
		.sram_avalon_sram_slave_readdatavalid                         (mm_interconnect_0_sram_avalon_sram_slave_readdatavalid),                      //                                                   .readdatavalid
		.sysid_qsys_control_slave_address                             (mm_interconnect_0_sysid_qsys_control_slave_address),                          //                           sysid_qsys_control_slave.address
		.sysid_qsys_control_slave_readdata                            (mm_interconnect_0_sysid_qsys_control_slave_readdata),                         //                                                   .readdata
		.timer_s1_address                                             (mm_interconnect_0_timer_s1_address),                                          //                                           timer_s1.address
		.timer_s1_write                                               (mm_interconnect_0_timer_s1_write),                                            //                                                   .write
		.timer_s1_readdata                                            (mm_interconnect_0_timer_s1_readdata),                                         //                                                   .readdata
		.timer_s1_writedata                                           (mm_interconnect_0_timer_s1_writedata),                                        //                                                   .writedata
		.timer_s1_chipselect                                          (mm_interconnect_0_timer_s1_chipselect),                                       //                                                   .chipselect
		.video_pixel_buffer_dma_avalon_control_slave_address          (mm_interconnect_0_video_pixel_buffer_dma_avalon_control_slave_address),       //        video_pixel_buffer_dma_avalon_control_slave.address
		.video_pixel_buffer_dma_avalon_control_slave_write            (mm_interconnect_0_video_pixel_buffer_dma_avalon_control_slave_write),         //                                                   .write
		.video_pixel_buffer_dma_avalon_control_slave_read             (mm_interconnect_0_video_pixel_buffer_dma_avalon_control_slave_read),          //                                                   .read
		.video_pixel_buffer_dma_avalon_control_slave_readdata         (mm_interconnect_0_video_pixel_buffer_dma_avalon_control_slave_readdata),      //                                                   .readdata
		.video_pixel_buffer_dma_avalon_control_slave_writedata        (mm_interconnect_0_video_pixel_buffer_dma_avalon_control_slave_writedata),     //                                                   .writedata
		.video_pixel_buffer_dma_avalon_control_slave_byteenable       (mm_interconnect_0_video_pixel_buffer_dma_avalon_control_slave_byteenable)     //                                                   .byteenable
	);

	Core_irq_mapper irq_mapper (
		.clk           (sys_sdram_pll_sys_clk_clk),          //       clk.clk
		.reset         (rst_controller_002_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),           // receiver0.irq
		.receiver1_irq (irq_mapper_receiver1_irq),           // receiver1.irq
		.receiver2_irq (irq_mapper_receiver2_irq),           // receiver2.irq
		.receiver3_irq (irq_mapper_receiver3_irq),           // receiver3.irq
		.sender_irq    (nios2_cpu_irq_irq)                   //    sender.irq
	);

	altera_irq_clock_crosser #(
		.IRQ_WIDTH (1)
	) irq_synchronizer (
		.receiver_clk   (clock_bridge_out_clk_clk),           //       receiver_clk.clk
		.sender_clk     (sys_sdram_pll_sys_clk_clk),          //         sender_clk.clk
		.receiver_reset (rst_controller_reset_out_reset),     // receiver_clk_reset.reset
		.sender_reset   (rst_controller_002_reset_out_reset), //   sender_clk_reset.reset
		.receiver_irq   (irq_synchronizer_receiver_irq),      //           receiver.irq
		.sender_irq     (irq_mapper_receiver0_irq)            //             sender.irq
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (3),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_reset_n),                      // reset_in0.reset
		.reset_in1      (nios2_cpu_debug_reset_request_reset), // reset_in1.reset
		.reset_in2      (audio_pll_reset_source_reset),        // reset_in2.reset
		.clk            (clock_bridge_out_clk_clk),            //       clk.clk
		.reset_out      (rst_controller_reset_out_reset),      // reset_out.reset
		.reset_req      (),                                    // (terminated)
		.reset_req_in0  (1'b0),                                // (terminated)
		.reset_req_in1  (1'b0),                                // (terminated)
		.reset_req_in2  (1'b0),                                // (terminated)
		.reset_in3      (1'b0),                                // (terminated)
		.reset_req_in3  (1'b0),                                // (terminated)
		.reset_in4      (1'b0),                                // (terminated)
		.reset_req_in4  (1'b0),                                // (terminated)
		.reset_in5      (1'b0),                                // (terminated)
		.reset_req_in5  (1'b0),                                // (terminated)
		.reset_in6      (1'b0),                                // (terminated)
		.reset_req_in6  (1'b0),                                // (terminated)
		.reset_in7      (1'b0),                                // (terminated)
		.reset_req_in7  (1'b0),                                // (terminated)
		.reset_in8      (1'b0),                                // (terminated)
		.reset_req_in8  (1'b0),                                // (terminated)
		.reset_in9      (1'b0),                                // (terminated)
		.reset_req_in9  (1'b0),                                // (terminated)
		.reset_in10     (1'b0),                                // (terminated)
		.reset_req_in10 (1'b0),                                // (terminated)
		.reset_in11     (1'b0),                                // (terminated)
		.reset_req_in11 (1'b0),                                // (terminated)
		.reset_in12     (1'b0),                                // (terminated)
		.reset_req_in12 (1'b0),                                // (terminated)
		.reset_in13     (1'b0),                                // (terminated)
		.reset_req_in13 (1'b0),                                // (terminated)
		.reset_in14     (1'b0),                                // (terminated)
		.reset_req_in14 (1'b0),                                // (terminated)
		.reset_in15     (1'b0),                                // (terminated)
		.reset_req_in15 (1'b0)                                 // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_001 (
		.reset_in0      (~reset_reset_n),                     // reset_in0.reset
		.clk            (clk_clk),                            //       clk.clk
		.reset_out      (rst_controller_001_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (3),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_002 (
		.reset_in0      (~reset_reset_n),                         // reset_in0.reset
		.reset_in1      (nios2_cpu_debug_reset_request_reset),    // reset_in1.reset
		.reset_in2      (sys_sdram_pll_reset_source_reset),       // reset_in2.reset
		.clk            (sys_sdram_pll_sys_clk_clk),              //       clk.clk
		.reset_out      (rst_controller_002_reset_out_reset),     // reset_out.reset
		.reset_req      (rst_controller_002_reset_out_reset_req), //          .reset_req
		.reset_req_in0  (1'b0),                                   // (terminated)
		.reset_req_in1  (1'b0),                                   // (terminated)
		.reset_req_in2  (1'b0),                                   // (terminated)
		.reset_in3      (1'b0),                                   // (terminated)
		.reset_req_in3  (1'b0),                                   // (terminated)
		.reset_in4      (1'b0),                                   // (terminated)
		.reset_req_in4  (1'b0),                                   // (terminated)
		.reset_in5      (1'b0),                                   // (terminated)
		.reset_req_in5  (1'b0),                                   // (terminated)
		.reset_in6      (1'b0),                                   // (terminated)
		.reset_req_in6  (1'b0),                                   // (terminated)
		.reset_in7      (1'b0),                                   // (terminated)
		.reset_req_in7  (1'b0),                                   // (terminated)
		.reset_in8      (1'b0),                                   // (terminated)
		.reset_req_in8  (1'b0),                                   // (terminated)
		.reset_in9      (1'b0),                                   // (terminated)
		.reset_req_in9  (1'b0),                                   // (terminated)
		.reset_in10     (1'b0),                                   // (terminated)
		.reset_req_in10 (1'b0),                                   // (terminated)
		.reset_in11     (1'b0),                                   // (terminated)
		.reset_req_in11 (1'b0),                                   // (terminated)
		.reset_in12     (1'b0),                                   // (terminated)
		.reset_req_in12 (1'b0),                                   // (terminated)
		.reset_in13     (1'b0),                                   // (terminated)
		.reset_req_in13 (1'b0),                                   // (terminated)
		.reset_in14     (1'b0),                                   // (terminated)
		.reset_req_in14 (1'b0),                                   // (terminated)
		.reset_in15     (1'b0),                                   // (terminated)
		.reset_req_in15 (1'b0)                                    // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_003 (
		.reset_in0      (~reset_reset_n),                     // reset_in0.reset
		.clk            (clk_0_clk),                          //       clk.clk
		.reset_out      (rst_controller_003_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_004 (
		.reset_in0      (~reset_reset_n),                      // reset_in0.reset
		.reset_in1      (nios2_cpu_debug_reset_request_reset), // reset_in1.reset
		.clk            (sys_sdram_pll_sys_clk_clk),           //       clk.clk
		.reset_out      (rst_controller_004_reset_out_reset),  // reset_out.reset
		.reset_req      (),                                    // (terminated)
		.reset_req_in0  (1'b0),                                // (terminated)
		.reset_req_in1  (1'b0),                                // (terminated)
		.reset_in2      (1'b0),                                // (terminated)
		.reset_req_in2  (1'b0),                                // (terminated)
		.reset_in3      (1'b0),                                // (terminated)
		.reset_req_in3  (1'b0),                                // (terminated)
		.reset_in4      (1'b0),                                // (terminated)
		.reset_req_in4  (1'b0),                                // (terminated)
		.reset_in5      (1'b0),                                // (terminated)
		.reset_req_in5  (1'b0),                                // (terminated)
		.reset_in6      (1'b0),                                // (terminated)
		.reset_req_in6  (1'b0),                                // (terminated)
		.reset_in7      (1'b0),                                // (terminated)
		.reset_req_in7  (1'b0),                                // (terminated)
		.reset_in8      (1'b0),                                // (terminated)
		.reset_req_in8  (1'b0),                                // (terminated)
		.reset_in9      (1'b0),                                // (terminated)
		.reset_req_in9  (1'b0),                                // (terminated)
		.reset_in10     (1'b0),                                // (terminated)
		.reset_req_in10 (1'b0),                                // (terminated)
		.reset_in11     (1'b0),                                // (terminated)
		.reset_req_in11 (1'b0),                                // (terminated)
		.reset_in12     (1'b0),                                // (terminated)
		.reset_req_in12 (1'b0),                                // (terminated)
		.reset_in13     (1'b0),                                // (terminated)
		.reset_req_in13 (1'b0),                                // (terminated)
		.reset_in14     (1'b0),                                // (terminated)
		.reset_req_in14 (1'b0),                                // (terminated)
		.reset_in15     (1'b0),                                // (terminated)
		.reset_req_in15 (1'b0)                                 // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_005 (
		.reset_in0      (nios2_cpu_debug_reset_request_reset), // reset_in0.reset
		.reset_in1      (sys_sdram_pll_reset_source_reset),    // reset_in1.reset
		.clk            (sys_sdram_pll_sys_clk_clk),           //       clk.clk
		.reset_out      (rst_controller_005_reset_out_reset),  // reset_out.reset
		.reset_req      (),                                    // (terminated)
		.reset_req_in0  (1'b0),                                // (terminated)
		.reset_req_in1  (1'b0),                                // (terminated)
		.reset_in2      (1'b0),                                // (terminated)
		.reset_req_in2  (1'b0),                                // (terminated)
		.reset_in3      (1'b0),                                // (terminated)
		.reset_req_in3  (1'b0),                                // (terminated)
		.reset_in4      (1'b0),                                // (terminated)
		.reset_req_in4  (1'b0),                                // (terminated)
		.reset_in5      (1'b0),                                // (terminated)
		.reset_req_in5  (1'b0),                                // (terminated)
		.reset_in6      (1'b0),                                // (terminated)
		.reset_req_in6  (1'b0),                                // (terminated)
		.reset_in7      (1'b0),                                // (terminated)
		.reset_req_in7  (1'b0),                                // (terminated)
		.reset_in8      (1'b0),                                // (terminated)
		.reset_req_in8  (1'b0),                                // (terminated)
		.reset_in9      (1'b0),                                // (terminated)
		.reset_req_in9  (1'b0),                                // (terminated)
		.reset_in10     (1'b0),                                // (terminated)
		.reset_req_in10 (1'b0),                                // (terminated)
		.reset_in11     (1'b0),                                // (terminated)
		.reset_req_in11 (1'b0),                                // (terminated)
		.reset_in12     (1'b0),                                // (terminated)
		.reset_req_in12 (1'b0),                                // (terminated)
		.reset_in13     (1'b0),                                // (terminated)
		.reset_req_in13 (1'b0),                                // (terminated)
		.reset_in14     (1'b0),                                // (terminated)
		.reset_req_in14 (1'b0),                                // (terminated)
		.reset_in15     (1'b0),                                // (terminated)
		.reset_req_in15 (1'b0)                                 // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_006 (
		.reset_in0      (video_pll_reset_source_reset),       // reset_in0.reset
		.clk            (video_pll_lcd_clk_clk),              //       clk.clk
		.reset_out      (rst_controller_006_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_007 (
		.reset_in0      (~reset_reset_n),                     // reset_in0.reset
		.reset_in1      (video_pll_reset_source_reset),       // reset_in1.reset
		.clk            (video_pll_lcd_clk_clk),              //       clk.clk
		.reset_out      (rst_controller_007_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

endmodule
