��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%�����d^S$�0���<SG���0}�q�hS���.o�o�X{R�?9�x��ּ�@�����Y�v.'1t��>�1M=�\,�i�R5V[d�M35��c��HT���"��3�xE�'o�wu����	UL�F����K���hb~˟�Oa�3:��mm*�{���H�;(�=��Զ,UH�X�����쎭;n9�hp������ ��u���B$r�䅚���I��+",��X��@$@���L@����rVj����C����4� �ҭ:�r)�1��L�
p����{�_��Ç ��g(/����@��Ȅ�J���5�.�*z"�5,h�A�	y���l�-��X}��Rq`~�ĽjB�M���$ń+>Ĵ!��Ե��8�2r�V3�t�ܧ��Ey�SL�ˣ;#�
���O���7U)� �ꫢ�f�8�5h���f�Ph?"ۍm�X��N�����c�� �<��`��2e��,G�@�wÏk�i�F8C7z�����j�0-�B.�}�(�h���+7��/�1�)��>e� f�Y�1�� ͞D.O�>L����2��Hm�pE�U��-S�Z����E�߼�iF���h�K϶�;]����,Z���tNW��W�v�	_�|�DBӸ�w����}$��X(q�yPo��6�NS�h�p<���L�j��5<��R�V���{ҪK8�t�=�1��QB$}ʆWI7�fL��r;K�Gd���."�P�R�����ȜZ^ ԗ���O$��L�/y��☌HZ�����=b��W�|������¾u�ǎQ�ϰ��q͒l���T��Ը4	|)C�B�P�4�u�	�7JFz�Ü���Q��|�'��:�/��~���K��>�+E��n;b�*�I0���+�EJG��R5�����J���n%����Y	�O�\��E�7H���Pɴ�sb=��������v�2 ���$?��:�i2}/�l��߰X�ZP��7����yF�,�t���zu�XQ�-} s�Q���C}�ƍ��0�̓�fT>AE��k	{�t^���~���v�m�cI1����ك�:djҥ��M�/PIS��	��9^q��vi۵f��Ս��ZS�KR55�7@�fC���ޓ�Ю��"Q:�EW~�Ƈ�1�e�$f��M���M��	��.����M bL#�KA���Ǆ�P�?I2i������i���A�f���BU��� \V���d�N o��hF:�#1���o�H.y����I�Uyb�c}��_��pښ�R��VᏫl��Zqz0�
�)ZI+[��$�M���Q��Lr����g��i����<ylkN�v��3�PH�[̦=�qAް��籘X�E���2���;�hQ+		.�[�!ˆg:WF�m��� d0UG7W�/�(C�!��xm:�$YV��W�&W�EC��
Ux���JQ�>����MtA�����C��< 9�L᠒N�/̲w��֩{�4ڢ˅$Ho
F���"�qэL5��jǌ���x���B��m��#�df�_��`]c���1�I R�T�B.�����x:.��9Q��E}�W�j�1����/��4n�{�Wܓb�Ԧ��X��¤k����y|�u��]�c_���_ʥ0
��Sٟ��$:��GS��ҳ����KD��?��\����W,�J��2(VHY�x��bbQ.�I���wДi-��8�A.� ���i3�P�P}�m���b��S�>o�7��"dM�JWP��c�:q��wn�fV6L�x���꣱�p�W�-�	�0���H����ë�|,d�|=�7'������U%hA<n�,��N�/6G1Pu��֖���_���qo$���~���u�,_g`H,j��y��!w�̻��!ۄ|"c���'�eF��4��[|�^����o 9V�>�u2\(i 7��~�#"�2�=�׿���q�꘵^G���f�Mz��=������M�!ڂEh��^#X���פ1-=*Y_�Ј)�E��8�F�ZQ�--����%mc2�������^��4vA�!�0`��5j�<���_n�UϏUicAYA��G��dyGzt�c+{0Z��=a޷Ǽe ZBQD����-��+�OP�į�T�^3BN�G�P|.)?��^��|o�XUY�9���1
ı$<֓��K�S�='�EˍO`�OquL�j��o���)o��e/;��q�鍼pUOe¡�H�KI&�4��R���{h�K��+Β�Xytv�b��%^U|5��&�=�WC��UĲWF']!{����S^��'�1`�_k믿un2ޑ	
��χ���54���pz����uc�\�A����A9��ծߨ�d��l����p?Td!�р���C�����*�]j�8���Ĭҡ� b�=��e3�[�ndH n�y��,�@mqz�j����`0��d��f���	VY�O������,]�Bl������2�B�f����^߯5��;h���e�����<-�Pg�]�u���x�0����	�#�iUз�yjg{�X���;j�H��a�r�_��<K��u0X��D`}rN펰2΃���T���0�08K��րZ`:�.\��<��B�!���~��p���㢏=�<'�W9;w8�X��_X�3!��F:��ݴ:,'���BI �q kL��/���Y%�פ��`��S��6=i�bh�g2y?�ւkJ@�ك8}�: Y��G�#-j#��;�o�YMZ�B��p�����R��z$R9��Yð�R-߻5�v�|�D�s�0�"i����4}Wq:=�cD=��6�9P�jHa�J;��� �� ��q�L`����ԛ8�w��|R,�sjuWړ)%:�f��s�2��d��X߿8�lw�����~M�$o-�P��{<���v�R�$+G�v��=���n,��kv�d]�<)i���Y3d.%ajK%�o��}F�P%��y�G��	zW��U����vwg`ᕣ��"�G�/">]�)~����)��]zr�<�d�Ȼ�w����&	y�c�	Fd�7��z��S�:2rښX�/�2t����Jb�e^��L5��yl�q->��:�c����e@��	H�o��40�/�x��4㤐Z�?Ձ��!���'V��'�:o���
�r��1��%��y��LT���0���_���^֎�JDj/�N�M����P˕������q��`v?3�"j3���	!T"���W_��	7՝�&n!4Rxi��H�ςʈ�,C冫�f�s}^��6*),���J[мR���=���ܙ%�1ᘿ�����a>K���2��y�(��]��q��V�?�U�,_�.UZ8'�C�i�Ol1xǹ�	&�C�Vu�%]�ٚ\3��W�C�@�q���x�� }Xj�2��ٕf��b}�c�僬�	;�~=)�U-�4S���a��'���mniyQ���FՈ�`!<d�4��̇�
p����;k���QI52��V��֑<'PP����# T`���;/o� @��sh'���.�KR���(���JW=a���HR�
 �;�bH���Z��Pa�̐k�1�(�$�6�t��+���v]��=2-�`w����[���^���>� (x�B���3	�5�󿖞�eSb1R�7�r½n��ip�l��mt�*Q����0~@e�fퟳ��: �Qg�	�y��l#s-ݱ\:�"��ώ�
�BjB]�Z�ZXlT����),Bnԋ���w�OM�4Ym���x3����P+}��OZ��9����8q
M��bܦ*�;*��|�8����W4-� ����~�,龓*<�?:�f��Q�Unq�~��� �&Bi9#l��d/V�`ա��M袔�n�2%��DJޫ�:p�*�`�$,7W��Ȃ�=����0���(��
C6U����@��C�e[\��1$�:�A{k�s=��=V(�zԴ4���4Y�S���P��rFSz䳸zpל�pŅI�����6���#����pVb[4�n3��e���P)� u��{<[�.���Cۖ����G.'�"�����˛��A~B�tA��+������1$����m���
�k��4MJ�҆"�Q�J�"��f/`w�2��I�0�r���k�:�M���zK� ���܈KFEI��x�K����g�_hU�\r�o�2\�u��SjO*m`���h����yK���v8��R%e�gR�J�1�ų!iU��֧#�[������b���}ϑY�����JG�|�]7a��.����˨�G�*����?_�tm�-��`��2�L� ~�T��DIw|e��7o�K�)����]��c�9*{����m��0���9'��=�h"��1sI>�$?6ݗ_ȓ]_B�^P��?�&|ʫ�fُVa��D���ai���IT@���c�"����A98���B���S�|}���JE���U|T9ǭ����#��賭��H�0����k�ʽ�=a�F"��>'$m�Y��P�)��J)cX�<:�_�&ѥ���A�}�/�/���z��+#�dp��G/����`�{�rOh7�	�YK�IV��*${	�8���?�d΄�3`�k$�/�.����ص�܊�2��������g��v�v�:JJ����Snx}4�3��
Հ��=kM��`<�����d�mF���Łr�����K�u���a2�*;xa{�ơL�nZ����oZˍ���~e�N>��ǔ���"�
b���<$C�)e���R����c {��
+�^ۦxL��ӝf��}�,FgU�9���t�bެ�GHp�O����|����Y��w��F���t6���=f���omPN��Ғ߳d*� j�ƴ�B��ҵ�sV���驔�~�Co��R�[8vV))�=J/Q��.Bȁ&b�̌�ƸJ�o-�+)A�U�F%6������t����:Q��1ږO�G۴�.b.�Kz�,��d�q��X?u���[�U;6/w�<�۫�Z��؎:��v51Tv�a�=$������s��}��8;�+��� ғ�7��%�|�O+�$"m	�?l���$x��O�/�U]��Ie���T�m�b]R�L�)p���`��\�ҟ��~;�s�'`m^$�O���h��-��oy `��������f<��G��⼀
ӜyBג�L���9��B�IZ�D+��K���ɂi��[���Qv���+m����D?�2y�{���@��_m��C+�r���Fe��ǅ�[�T�_���cF_^��5�)y�� ��ؤE3�D$2�р�sl�yw�M�aP#��渆�87�W�˹�f��{���\��Ǿޤ��A'x����L��sVM�rC`�0�)Ei���S�xi
p
�d9G��M[�I#�-�� gl��� bC=-�����i�*����A�P^�m�*fi����d��C,$Q��r�d��#.�'���&HV��F��@��o�����!/Bw����&`���H
K�-@�P&����92����D��<J����Q$~�kI6i����&#�S�ot��<������c�%�֒��c��18�z�ϫZgs�܅����\���9|��I=��s�����"�H��Ϡ�v/
<B�x��p��^����?�-��)d�_��=0�/�����ld��>�˺��P�
�O0�ca��B, ��5*`."$��7,�u���*��d�>G�h�K�_��M��COr,�|G�*x�h�Uy���xOE���Vª%�X���C7Ƃ[s;���j���+!��n�t�o������.�8�,ݧ^�0Eas��c<��
���b�}���܃F�R�"�'�?^*��.�Z�|7uC�jBhrC�"{,`c�-g���خ�6�kY���@�@Ahs��.�7����-[��8�,K�#%ӖБƘ-p���Yi����(�_7���je��l�fmR�?#�5��C)Ũى���4y����,j}rŰ�☉�Ô?.q�z�LV�[�ǌ��>;��ЍX��:���k�CRY
وt��>v����|'@��^�B��8K^���q��gd��/�?����q���ʎ��Fr�K�'߬<�G�Sr�<��b�Ƌ��4D���6Q�7'<�1N�uӵ��b�Q��?�n���Cŗm��.��8uy��kZNF�B���Fy��H�%;A"+�s�M�X��j���o���E!��x�3Q��&T�}tt��7���+4�����������^�G��og@QA���H��Y��F��vi��3 V�q���9hJ[�.�I$�GA)RM�6��װ�P�k���|�gǈ�)����^�a��DAa��#}���ۯn�sjc�E'9v�����k�X�	��9�}�r;bSrX��oF��~!��@�e��w�����n&J��F������L
�t�5�BZ����=��<���g4�;�1����hm�p�7gF��AŅ��d��������q�a����+I-�w*>o��Sg�L~���c$�̊},�g�y�t�/��(m�9�GchG�m�+{�F�J,a!JA�t�uG�0�ܠ(PA�`��S���\a�&lr�D8@�ڛ��������^��;ϫ(&��w�o��tĂKB��5z��ІX��4n�84-mO���x�>���8���Za�D��z���)�y�E!��a;D�,c������Jnxr\��=1�x�ױ8�z�I��:�A\^
b�
$PX$�U�W���<}���+��@@�u�0�c�v�X���%���L�C�)���=�_K�
���YU�5���0�����Y��h-05Ѱ�� lH�U�}�׸#���;SC��k] φ��)��A)�D��cԋC�E���\�X�?Zu��3�s�7_�`|�;����Q|��E�D�����5@��P`E��X�,��L�F�8���p-��*	t=��{M`$���ky��1��QUx���\����m�?_Rq��H�[ĩs.��C7�h�`�URe�E�B�7X��E9��O�Y�`,�t��R���jX��[O�td��;�R�oX�wQɿ����?��W�XWs��D��k��������' ��h��)6K���m�{�j�4>��#���E4��K���q�cBW��}��r��ĜQq��'�ȧ஻��FW.���B�B4,TUQ��Ɇf�,M(d��3���wx�^��������_O�s��}⒖�,���f\�&߮v�X�_�6.�t[�aEVd�I���1n��{5�ڤs���AoU
���n�i�KU2%9��'���Y����
	ŭ����vW��]�أ�W9���sT�� ��л�G��� ��O����n���U�-�Q���u�|��0vt�<W2;��� '���Gf_�~A�ΧE��}^�bw�Uw��ʰ���w�r�J�a��l}����晶 �:oq,�#�I��OD�v,3o.
�����n�yҩ[��ٖ��W�%9V�cY�%�F|�d�a�0!���C��z�X��tr��������U*!�x�Jj�����Ny+��OMyB��
�TzS��;��]֡��kЬQP����:�P�&k٠��BM�5ܼI���~�Y�1]��+v1�
4v:�~N�/�e7ٲg>`��)6�I���ÊMb'1�w<�%u~��~���]S��ǕC\I��1T����'<2��BM��9�vvQ|���~�ߴ+� K�o����˯���ʁp=�� zO�����]�k����Bd[ 0Hj���z���-]���|!.�"VX�66��,;�	X��09��L��8;"���^A��̅�`~��F�;�M��x+�D PjϨ	�`';)c��b����dC��U���]4ש���rĸF�d�
��&�
!/Q���ā Lw(4&�p'ȵǧ�8ƍ�4W+kmY@���P��oԨh�*O���Z�g&���'�^�{��s/³�l�u�Ǳy}7�Ű{=��)�ZjnA���d^J��
N�Es�?┥�AJ�[��J�L���<��J
=g������z��;����C���	��J�Щk�u�5�K5�\=��v����`/�8s;�N6�(���V j�@@��v�y���$U��}�o���A��4��ښ��ƨ9@�����Њ�7I����<�@HrS��o�v�vg=.$Z���^�I47�J�Mia��D�Ǣ0/���'��x&� ��2�w_���G3���tk�hhX�~~�#�~��Vk}�8����)� �گ�s�f�s�������[:��O��@Bz���������7�3/^�����p��\>g���#�
E���f!����E��*ΨT*q���[ܴ��M��F[��Ų�H�cG����t�삆��Z��ǀ�b=yv���{�%��m�2��������m����ߒ|�1d�x���>�K���x���8&M�� ��i #B`���5����N�]�7�NQ����{|a�Jl���zFƑ�
��IF4�>tOKs���K�Y���Z�5�/�N��A�"���Qz��z܆����p���l�d�{&h��j@k����Ts^��������D�����j��.4�cG��(!�����~'�Iyq¤A�vjҹ��7��@�v�@��
�B�\����d��"�t�j�
a0<�>���P� ��a�"5�z���sݛm��X�=���s�h��M���)���D�t�
z��l �Bq�������e��2�=�WJ��_��^V.�P�y@����p��S�woô�bQ����?{�a��O뾂d���?N~׬G|(n�<�fHhy.�v�����3��x�SAh[���*�x�-��+@�e[�-P�� Ґj���0{׶�O����IL((�_�y��b��a7hoSkBb<:ƿ������ ��[`W;�b�	-�+bM"��\u�8�ߒ+cs�_@9�d�Z���Մ��z?�ι(��Ϙ�,H�����3o^�vO	Yp��v��v2.�Q�~� B"�$I"{m�%g�`����n�� ���I�Z�,�Α��FT ���βb&�Eƿ�9H��� `��msa�y�+J(I�N������to���U�Q�[A����KG�lV�B�}9�5�����v����8$,���OCӳ]��)��N����j{Gy�&J��x���]����
5�C�L%�b��F��м�"�?��'] �
��_7�_�o;�] �°��6�8uv�P���>��� �a�I>m�*.с��Ɖyc�LXU��� �:�D�"��ci~}���>tB�%E�b
�Z�z»�9�@\t)��4�/0�T�&VW1oFc�[-���[����8����M8��Gh����+�H<�	Wi^�6-��[m�o����d�+��'�y��)������b��m��0s���VoIu��%~l�DhSZ{�&�z��M�r�	���h(����y�*d::�l�{�@�W.��EF���8�B��7)�8�����O-O����J�Yn���u��gN�L��s} >�r�@�v�ZH|s���q�o�����T�Wim$4|�8{pA{Xz&���@!#|�_W�"B5pX�Zw�3��(e�d�h����#c�7��?ƙ�vjlc��=����lG�=	G�ãd��QY��>�б��~	��DK*[� �e�r�ؖ��d�UNSU%���"C��P�f��mBW�%��1.#��;o�"֤��'��G	�
-��u��&�B�J������#���Y8�h�{�G��~�S8���ӿ�������mdA���m�Qw������U�
�C�&|��"�э]�*��ץg��V�Wjb�&\�hS��MD��!��:Bs��gLO�K���Ԇ$DG�#����I���Րԃ�&©AA*�?d��5O�xɉ���)�IѺ�l�	��2��N�[��zB�ş�����|�ic���i�G�I^���L����ѿ���uL`��9a��B(?�_�\��D4�u"L��� >���գh��7����e		���ץ=�B+���Pd����ޛrkh�K�Pt���M�Y���ʯ��W�`l��'����z���û�Rl�t�J�O�uo�#�������~fpZ����>L{.	,QoX�z{��P��a{��4	-����ݩ��v[��g���+��
 ��OZO;�܂S����k#"��~�U+�q�����[��I��� >-�g8(���B3V��pڡF��w��>Ո���hM-��o<������O�1t9����
(l�l�:�	1�$�ln*+Ik����~;�C`;�M.Cvq�๮aW\���B���'2<X�a�[*�����(?A���-������K��׃H����/�oę�ǔ�i����b03�צ�ىZy&����Cu�_6��9q��Qx�w��r��Rn�俱UG��B+mx�	Ef2��d��x�,Vzk������Ma�1q)�\-�W���&�kh���2 H|@OIK2<�qm�}-��U���B��b@�⺀1�|���MB��VW�A�5���>�q���'������͊�N���z�� j �2S���Q`~�PX��(f�#�=)�����-q�{���
y
�J��dF�!��(kɊ��Cx�o��+k�v��ax��ÌB�=z�t|{-a��3�X}��"P��s��{v��w��XX��3��$}�"���F_��#~B�z�Q�,D�>͋WY�y�HK���^�o&/�#<jd�f��"ԅe['���7�#Rӎ�#����oC�(�|�	�L����Q!��]5���3��4�����.,�A��8v�=�庎�(�[�f�ҭ���:�����c,��l�>��>P�;�����[���"UF�d��濝���G�P3�8+�~�
�(����s|��M7F�悶~{Jf�b]]N�caJ^�En������u�r��jE���Y���I�0��:zt���a=�	���L��$A�-��M�}�k���*(\F���m!��k�[�G��RU@$���D����M�/����;�����x$�d�z��И�yZwj?��r~�Y�Q�;l�F���)����? ,�ׄW4�U���a1Б�RW�ʯ⃉
��j8���*��/Y�/�$�aIڕ��lY�x�O�\�Ù �9*Jܨ�	�ݻ��r̕�D~���D-����=g�>Ds���d�^2C��h��ɱ������[���odRv�"�zЦ:)'f���&�Z��9H8X!����
��[o��>�����sG|�.��$ֿ8�>+dJ����{�4���H+��/Z����nC�?��7�T˦�đ����A�c�e�rF:�;˱�V@��慇��}�8�d��Gl����LI���a�q�5�vڱ;@Q_(�$��/O��~�b��?1�����	��ٺ��	�{�1��y���	ف$��c*j5��Z����gW���M��Y��[>����^#S�eP*�7i*Q&d�ћ��`�v�T{��8���6ޏ�熘���x��Q�T�8�J�W�.Ʉ�
\8�}���|�]�ɽGc~W R���F)��j��	�&�P�a5GK_�/6	���t�JEY�t���p�
3��s��ھ�g��M �c�l, +X�{�F�Q�Ȫ,�q��k�ӂ��Br���{;؃T�N�A��F�yo�~9y2��U7��^V���6�h�Ƃ'�ß6��]�B�,��i��=j��[��A~��?#�A�A������޺����8�k�e���`�lB�x���9��nTl�2J�����B���vXO|#l ���� ���Ȱ��A$v��R�t3z dpUZ���}2Y���6�~`�
�|5��$�v�b:c��d�6�����&Q�ב�#�
wu4��[5�������6�������GV��#�X�x��>%p��/���Qh洪d� ����4MڱVG�h��~�-0�Wr�#=rE�r2W�
b�X@�>���WRRмfH��2�/P|DU��`sPx��|K�um�����v�D��*��)M/XN�YƋHa8�s�7m�k$mӈ�-�YX(���������}T}�ڧ���pxW���x����/x��T��%䌽���)��O4����W�Z�{U���P ��uP�����������8b�L�p�֛�݇#]� 5�����ۓ�E�x���?}MU����t	_<-����c�q�F�ܶQ�_��'D,��$�'���!����疳���� *�Q�s����<0n,/��T�K�s�C�(�7�~�N֡��C6HЂ"���|��/�ߣS��Z�?��~*@�I�$|��G��]n����c���8ږ6엧ނ�C!�������oň '�k}`�u����"�WI`qk��x��)�6qd�fr[��� �1�-�tl�xP��#���ٙ�ؐ�O�)<��@�I|R�r<�Yw���g�<�zR���X0���ǯ��Ƭ?��A�P�O
F|2� �Ҫx�g��78���;���$��%��.-E��9��1�M�l]ﺅj�mު6n�=��?���˱���aVwu~����N�02�-;	��tj�zC�X=�I�6�HI��5�ye��
P;�˼���n�F�V� bu>[���3�ʫ����!m��+�����7BW���[4��E��&�L�G���2��``w��[�7��,6D,���7���c]4��	>T������s��Z�w>nh�]�A��sd��1��1��I��ݶ�X7zx� T�k�8�����ƈ8�˧t��'���.V��&�W	��Q�m\��&��i!iłe��@ҁ�ʎd*��������_�~�_m�v�7X�Ij�O����yPNk�([*�]2�b0wB�uE�Z��J}�뇛�w��~X��Z>���m���r�ے��/W�h2t`����l���B5kDz�}dC����u�aK�v�/u-�Ϋ9�.I/�F��N����5ކ��7��"��v�Hބ�k��*}L�0�y�j8S�jt�ʷK^��E\��rޤ�\n��`^5zl(�����:Oɉr�DmEg�C���.]��&�x5�����>�Su@�h`E����Oݻ\���?��>}&gD��-95����BŌ����=S����� �����%�j��ft��m]^6�3jk�������;�b�2�dk�����
/)@���YHT�� :��7ɸA|�`h�TU������r��Q�`�c��qFGR���L��u�����T��a��;����/��t��Y.iĿAV�e]�R�_���$��$�bH1}�b�l8{^��'Z�}B����:��� �H���xU�_Ir�qBžc���u.mWX����ɧu6�X�ÆE�FN=�ơp��R�%�]�W��0�M<���sm&�j�)���r� ��sU�_�U��\o�պ!SW �;r�s���c"kȭK���E�����I�JL͍Q;��XN�q�n0��ƁMZF��a48e�ND�&07f8�ő�݇��ԲRW�I��5�����b�҉.��B��l���7�RL=�~R�ك���x�>��̈�(���UO�$e���� ��^u��V=�z��U�'9l0cU�|͐F�d�e ��E�p>-ƌ
���:��h��P:�l���1 omZK�NN�d����鱕6'��p�3��N8ms�}����vz�k�/p�O�FR<��=P8|�.Q�!��ɽ+�����;��& �3d��.�h�c����~a.����&�B��;��(7��T�>��	�C� yt�1Ͷ?��q��	��f�Gv��.Q�%�����i�/ޑ�sz��&<�p~,���)�X���=;�;��L�����w�=}��tp$5�AX��L�o�D�*�a�|���JĚOϥz)�ё4��s�Y���T&k�񥞥��{Fyw g!�X*����'u&���?��,�&�&�xL(���e���I�%�C�8�{�ɒ�Qx�IR�M;�r���S��>^G�*���wT	��A����C	,�-��P6��)����l�_�*�s���)��'m���*��O��6��\5�!2f�?��!�[,,&(?����(����P>D��@�g���0�B�1/����o[0�5���o�Ob��-_�9��T��D^Ø�BU�`���7b96��&w1�[ҋ�(C�%iپC}ʔr��3c�5�t��@S�8,l���)q��׼̚IQ�CY�E�<�>ĥ =��x.\�hf�{���Ơ�e��0n��J:�}��lV�<�
?�B��>�`���P[�(�>s�0����0:c.�fl(�~&��y.�I�K2�
0N�0������iM�c�wTdu�p:���H?#!-{�7TʐR��G��+׼��;��A2i.����/6���j;��h_$H	.�0��9zEPxv�N�*Z�jj�-�L[e���:���y~�c��s����i*�9UWj�ی�!B�D�)�k��wf���V}�f%Q��r-���KϨM�l�b�O���/ u��y��q��DuwU�[h�f�ac�ǂ���!�˝�x|�[�&�����%�h�v��[�v��?���5w$?׀Ԏ�ֿ{�bXאܓȐR��4���.����n�'��W�>��Y��&�tV^���K��QQ��-�|�{�j�����"���R	M�1���>�a�.|��2w0�+�3H�G�L�^��<
�N�$g�kx�sz­ξJ��D!cv�*�c����qS� �le�(iC	��)7RA�'v��=��ea�D�x���-��Ӻ���ȼ�h��껅f.�/�S��{@�,�x��xG��^�f�Aw,�H�cXg��}\s*�t(.]n
�!;�b�g�4��N;!����U\����v���Y��ꏛ\���q7H�c���^d޻�{��M)��a:g9w����<{�ZVS�k���ܘ�h)� ����Kl�y�՝2��2�rI���R?>�&��Ʉ�;�>���s(}��G�-]��;��@���:��#4�E$�@�dC�08��LS��P������Wy5(� z>h{�қ��R����K�˥ndy�e��Y�.̈́�1�C,�Ć��U^9�@ /?��y	D��Oc	�7�\��0]
Y������ET(�{!Ei�U�U�*�irx�-ui<(�6�^2������K�E2�-eL����e�}D���LI�hWX���?4�� ���j����4Sͺ&pN̙�W��]
q0.Fƿ�VM��z����F[2���DI��&P�(�Di��\�*��n�.Zb�NI�A��`|S�`�6wqQ�nx�@�K�=��M�P7;��Z�gY\s�h�"EQ�l*`���N|�&���2�="c�T	͸E#|*�z#��G�B)�v- z�n�@��;Ʊ�)ɀ��'e��,�����g)|MR$(}h������9��Sဪ9٪L*E{m�b�P��`p��:��̅]$�}ڄ��dD����O�e':v�TI���~+��t�t|�O���	��;m���.�:��ڬ���e�L�fb	�@YG%H��B�݁��m��v��0�" ȓ�W���(�Cq�g�n�C�Â���ܬ�s8����b��|�r8 ��	m�q�k@�!�r��~��?�ݼ:� }>���WT�/b<l�w�$ʗ���dР���&�����r�d���g�i�kbI�xc1���'�%Aq�n��z @�^���.������2'�q�z�9�.!���zQ%�b�O�����0	��z�DQ�K���@�F��m�s:=���a=�`�E�J�)�_,�A������������A���H��b���(C٥�ž�ey�������&���ݹy����HO����-�"��*�`>$$v�&�?G�ۮ�.l9��D 6wVP�Vj�T9�%�z�2x�#�*�B!y�o$[�LW�G�=}���������LUg)0y��Yaeo�~3
����/wn������U���� �-����r+�+#Yu_���Q�`[՜�f^BC�����Z�3�טY(QFh<�w�o����h�6nc��>�m� �Q$��Flad�)$Fs�(�AI��L����ح��&���^�h��� |��!X���/'� �� P��l܀1�z0�y�k3lMzG6<�Z=��HK^jD�;,�~X�� N��"�vFK[KO�����dу#S�#@�F���M8vh����,����d'E��:׋�f%J�]Ml_�GJu�aSթ�#��"Ղ^oBy��5e�I*��Y����K�n��p>��~I�o�+C��p����pI���V�L	�&K��%/��� �5�sv�el�L�ŉ�~���~T��� 1�jVh[v5���!dc�]y�K��p��z˧Pl\�H��(1/܇�g>Mh�eJ�U�[�3xfA�H: YV����j�c
d���uh�M�߻pCo�\���?` H���\V=H.a��B�Lg'��).���;.�O�Xm*8���3����N��K�����2����0�������E摩����C� �^�1Ϸ����e���Jd���0P�k�1U}��ޤ����r����~��7�&x�Y����&�b��D�Tb]�f�2��dij��,$�+��Q[q9�,����A��Q^Q���e*`���qa�4m&)؆��\�Q?�*�(m��a�P��v϶����Z�Di���w+��1F�w
�� �� �ɗj���h�WM@��8�^��!�s3��r+P�&�h��px��_��#l+@�x4| ],��/9��ӥ�
��J�YL�#E$A� ���D�����OHS|G���Өׯ��dF���p�^���-��o������~;aIZ�P�ᐦ���Ż�3�*�"k��U��,�1�BpT�Έx��~�*���:�z=�L�4��+q=W+B5Mz2A٫�����?���S�m�*�GE�O"���g�j��U�a�8V�Nv�e��$��ܰ�\���I"�R:H��6�����5��MD����D���!v��=�R�A��B��On��F���)P<�n��o�;��~
Y�t8T��~kt����?��;��<h���)D.=K�.�N��`5��Z7��.��3C#�$���X��*�C�H+��|IQ�+�%�.)���%�U<k�� �:ߌ`�zFqa�D\�����f�`��5@�7��)@x�xb�,څ�y�7C�.'D��r��S�:���)�K;X��5����	�.G��wŽ^�{0��R�,,��t���`�R���8yE����Ɵ���(�V�S��ʐo�g�a��6Wuj��4�:*��ֆ���9 ~cdEC`�~
��._)��%����B��_���w�oM=<*��N5|�yȯn~��ꬣãE<���	�FB���W��3�@Tr/\���J�'���9Q6
;����xm�����r�W)�� ��7�"Z}geJ�l�ՠ0�w�!��_o�y	; `�$���[����.1�{���#:ԡ�͉�D��?vEԘ�Y��?(� ����y��\���~�j�T!�����h�0�	S��q����!�mx5gq�U�y��*�qx��x���wB����g���0^s����C�ٖ�nm�z���'�O��X�����c$��(Y#�y�@��K�Zֱ)�W�[Rn��ʀ�N���s�����^w�̄�$do���[����B�SG�I�0��ޥd�P����j�H���o\S~B��[HrO��[���}V�a�ַ�{��c���f��T�.]��	1)�3Q h�p<c1�����S�j��օH�﵂8/K/UZ�Ed��X�[E�D7(�Qu����c���:6�|���29��,�%���kD'��Ƈ�ʿI̿/ ��;qل�C���E�@�u6 �{~c�&��p� ����wK���� �����C��n��(�e
��ϻ�P�R�lQ��˂\�[�=�S�ᓐfL!n�+�N�����9,�{�}+	i�ͣ/g�¢_}`���Ѹs�,_L�L�%%;�S\��"3�ݢUQ��ğ��B�\��r���'hF�$����qvod�LXeLH}�0�4��,�Nt��֞J��F[ڞT>��Q2B��B}�^�#�AM�x�@ڐP��:��u�Mi�&a>���o�����e_~�ibJ�:g��R�5t,z[�+@׷b�/#���!��Ud��R�_ὤe��1�(.������t7�5��[�IBz��B��lA�m�N��P�Pn�
�'��7���cz�B�qE/v�j���^�S;>T M1R�V?>	��_U�&�S��������I8:��D}�+/͝�,P�E�y�B��M�ĭ���Dt�h�ɭ5)��"kP���޲��Ǥp�5pQF�s�s�C��$g'�Q&6�8%n�p�gܾg��=�Y+"�i�z�0��r�k$�hn/]�u��S_��+�zh�UQ Na�嘠^.�M�7h6	*邇G��3E�,M}������ ���ַ.�������[ v������\V��:r'�?Ob=���C�o<���yU�^سa��I�j�;j�9�(�X�)3���2�a)�O��=��`�:w,|f�Q���7~V�?�L���J������䪌lna��61`��g$�B�4�g�ƶn����w�
���ڒ��y?�%��Z5�6�����j���RI6�j�u����lfh�><wxyR]�^�;���z �@�$F�LG��<�/���Ӭ��7�`�3�{�;��C�5��N�o[A�����yI6�W�u>N���J<$i�^Z�8�37��Ǟ}p�������2�,O����m~�XP�O��d��d�lG�BsVG������J����M
� 51���?�yX�����>�V0J-Y j8����D֦��9$u�&����336���A����gQ�W�֠����^��=����uW*�MFH����f�+j6�a	�y�&�&��d��h]�Ss������+o�D	�3�]�'��\���g�������|Yj>��bdQ�,�8o&|��sE�t�TKx���
mLF�bI�&��+��ɾ�Z���o�Dg���H�m'��H=�z���� m��!t���vy����/[u
�,1�ӣ}b��?�QS;�&0?1rU�K�Q絢Hf�mU,B�_h�<� ��Y�s���oTW��	�{=�-Qe�^D0�X��b�c�g'�����ĕ����vZw� ��"٢�Q�[Vd�(̪�����{)1V�z*�&pm����K���K1��<����k�<�P��<����<z�;7r�ǿec����$f��Z}=�5Y� �Qj���4�8��v�'��!�D� iʡd2���']��Z{�t��
m�*�7b4����L��/}�݊�Z����2ٺ<I�M3���7qhs9g����
�P��-]0����=5f���_�+�!��2��`�q�>J��^����ק��t�t��K���������$�\��[��ћn�7ƯBg��fv���z�X!��VQ!����.,Y���D+6qe��e=���1(J�z�d��N��h�	��dk*N�c�<bS��� ��]�,蒄���x���D<�zyy\^@}?��,bl��RUg3'�$��E=�HJ��Zb�*�c%��J��@2Ϙ�`5�����N����ȶg�#2-A2"r`ãT�����5��8]����V%��B���y�~��+���!M	Å>��`�A?�T�����<�q�2�"�;��}��/8�����K�ܼc�=e�h�1b@
��U�l��'ڈ�O��	���0(�y�oty�Z���r�T�|Ò̍�����9�µk��d�m=Đ��ֱ����CWe�����ɲ�:*�~�J��T�gR��ԙ~+��u�� �T;�-kjF���gD������z�Uj�4�Sy^���!�B)7v�ëO2dxy4RH�⍴Cȵ��Q28���m����f�ŭ�y�F����	�������$h��Ҩ��v�g���;ll�FYH[N�Itު�<L�@��������mn�z��fS�Txwj���r'�����Nm�YL��j`=my<{_O�`�HD����H�����
j�`d'f���hoCr{V��l�8[�[�?��pCtOpp��b��:�wS��y �ar����/�~3}\Kf���ȝCy.��e*�����g],5R�������;��+Y1+�F��mb��r�q�X4���k�>����W%��d^Iш7�}{3�42B��F�ôN7�P�}�o�yOafg.1G;����-�"~�
w�[)�tӺ�ԧ�ڠغK�(��ğ�f��؂+���T�<�%O�$]�R7�E�~*�Ƹ�(�"V�~�d�%1�� �}���lG����40�@���+�.ny~��R�.���[�d��.e�N�,X���I����	�i	mW1/G�?+������/���4K_��u��٢��]5�Փ�G\��|"��;��w�<Y�f�G���<?��m��B�D-���6��*�F�M�b[���~��2��H�&�`Ƙ?�Kk�c�w]��bTG���ƣl���Ϯ1�%\�ֻt�|aڶs-?$_�C�����V�l��6�0��6�uf0%�$�\F;����n[�4�0�:��x��\�ȥ}�f�r��:����bm���\�l\���G6�+���x�8�����=K?J���A�|��q~�:	�w�q!Fo򛘾�W#�'��M�s^4.���rd���d��ΒtI��Hَ�H�1DVک;m���:I���`gznIk�i�Ȇ�������~���Z-͝�I��j��uR1�$�=����н�Ė��^��7T�cݵ�2�����]8sP���7�����'����;H�G���X�,V��SN���|�j1v�F)�;�4j��{K?�~�f��c�w��m�gRWp��΋O�:9@�����1 ���A�G����B �aa���¶�ȼ�8�$��zn�2Ddh{rRE��e�ݯ,�q���678�_3����5D���B�2���@L@�d����Xڶ?�S3Hiz��z�����N��N�e��(H���x�լ�=��'s$0�>���a]D�@�q`�vO��7Co�ó@��4�A3�y�3Ҭ�ܓ�����+χ�'Irb2�2�DM���ͬ���a����[�<��ʰ��sv��b��=T>X���Yݷ�C�;8�3�*8��{|�d�ڭ9��
��C�.z��/J�C|��_���|�K����&\C��p�8�Y�Y��G�'"�^�k� u\���LT�
 X�.t?��`:�5&sY��L�[��/Ay�3^��'� �� {�o��4����:-�5��*������";ѶTFO�a�������P��}w���VP�E����;��-�#82��<����1	�q�\��blf��R6��?���B²e7�ET�#ٻ^b�|g�=���O0��ժ�Q�-�L���M�\x�>�����Dy�ʇ�8���+c�ǆ������{C�Q�,ʖ�L���+�2LI�T���08���mR�s:�$_�gŰn��o���N]��E�� �T��P3_
�������?�J���$������X���H���L1�4AS\��=4�)��Z�?J+O4���B&��2�M����ȓ��ZE �����;�ȏ�� ���d����ؾ�:ڵ�8��N՞��s�I��֖)F͛L7+c��Ā$P*B�3�Tҧ�|�"w>������T�� �Q+�5��$�%��P��e��6@EM(��^�w	!s�~��1�0��?�ro��;�\.\ǌT�x��(��1�+uk�w�✼Cq��m��o��9�U���6u�'��i���ŀn��<x�-�q��F�%nU�Շ
�#`>�D$/�m�X�P�s�[���)�q��;������8jI�E0A�`\���3vݽ��g裶˚��#5����1X)��](������e�A�Uz�e�C�s�t�����측��F�4e���x���t�,�t��'�g�>=܇Gn"���3��X+�y����˱��rS\�o�C�gC��޿�wZ�~�Ӳ}�#��1�\��-u�I�<�2���W���">"�2��S7Gl
�Ps��߂�pL����f.X�h	�fe䉻��}&;���ʩ>,N�T1R��t�>~�!�����A�C��y���}��5��Ws�?T\����5gZL;�k�r�ƒ]�@�&�y��{���K����,���I{�cA?��T9(�d����S�ԠM��7�}-Pp2Ft'�����E��q1����ޟ��*�:\�Z�|�c��Ζc��ȃ��$ｾ��e�G�&�U-����zښ�D�ɠӤ�F�W�b���vp2){�\Mn1�B�aɁ���8��(��Dz�#���`�}L����M��7W���_�#T��>s6�ߒ��.�/��[[�̓9c��Aᣦb:I�ҡP���/P�!9�&D��TvsV�4_����J���¼�R�[��?L��,��cY��c&K~�ݿ��;~��F�]���+���������3�fƬ�����A{���Hk�d�O���
���hέ�_q��7(�cSZW�<���4�?o�F_�]9�G\�5� eh�6 A�O���C����0Zk�D�k�d	wA½Ǥ��G}c��M�G~\b��h����~ٌ�|�U��B�'t-���g�p��i������F�
��bMf|'W������l��"z��I	�s��ړ��M5X'���6NF:��w�ؾǗ�@YD�� �%@j �0�p�ʅ�1�) ��I7l�3y�XY�����z�չc�'��]����)��&�����Y)��V��a�yz��7�H��TB��sY$X&ˮ��88�� ~�������m��:S#M�V-"��܁�}eV����'�8EJ�����$���r�6���,U)g�j��8\M/�;y	2��J��_�:�v�M�~����ҽ�|�=����]��T���g6\���U�� ����ԛ>M4�����FD0����掸�|h�)�~��������cZR�>�Mu=����0�*A�]|)�?��-2Q�%�.���j����sy �Y�1\���3VYAi	m�UZ��*�wYbW��k?�K\k��(�.�����00kX[ٱ:�Pq.fQ�e�Eهr]
�J��#���2�1�f�.0����t�=����$Ń�{�}ULRN���Rۭ��B����7 2�)L4���i$���?*/qo�R_��*5*�xu�YY��G.��� �J�`���B�J��nZ!��f�G΅0����3[C�� �\�i����v���l�|r����0���a�ʰY�D�4�I��0�g�+����f���N���/#��Z�믣�P�oS���ToG�0c�������E#��;����X8��0�&p�'T������%��E�q㰝��І����.F�5ai����2ϕOS|6.٢PL>��U?�ӝ���ta	�ܧf��=�/*��j�v��W����|hO��t@ᑀ9��^�N���Ť�/XX�Hǐ�|��ǌ+g�F3bTJs�~o���a���b��ɩ<�x�(75�kN4'&�6%;��/�O���t����h;��/Zf�qHu\]�"|� y�,��K�1�����+�Z1g�����/�w��,��o��W�^H˷�M�B�Se��T* 9�� P��9��K���S�>u��4��m� mN�0�m�T
��Y8�ұ02�=}�������,*a?�!Z���nC��Ć��"�$���v�l�+H>.�n*��P�-~!��	�Ø�Uz��"�bgs}I���17]U���V�$��.�E�EQo,��Q���� �oB��u^�AD��cynǚ�֯oS�5[zb�7b�&�$%5i܊�l]�T%�%����H��V��w)�I�`e]�5��`v����,'�c��*@��F:����^r������������m��AaK�In[.���FGzYj�3�aH8��ط�@�=R�<@��@"�=�9'TAe=|M*!Y�I�cs�W�<Y۞�$}`i���'���#��K�%���a �G'��H1�QZ�W�I�3@o�A�,-J��q���D1�y��]�P2 �=��z�6kJ�v`�b)��Q˗�)&�\<p���&}�)�9)�@4�f�n~���Q�K���+���a�<���𩃍O�XŇof4e-�����U�F���0�>�����e������i�71��z�èb�.�I�}6_�
� ػ���#�'��uY�ٶ٢��H��A�o6�4�T&]����'��j ��
���a�g���H�����vc�x�O*��p�0j���+b(-�����:]�����x�D���-^AFzO~��_s;���sF�!�{ϵ"/:}�.��i��~�m8�z�O-�̓���SH��GO{�*��e���0h	"uّ�n	��bg@���}���H	ge/S�Q���q�L��]���_��"������nƍa�4�_:j�.�5>#\\/	\n�<��Aa��i�W�8�	��,f��R���*[V�&zT���Q;q��&9t��gߒ���3.��_���@�h`��#o���-�:_�^b4N�{���j���}�g+���	}P,u�X���� ��i���E���N?VU�°�T[X;�l=�����[�L|�@L5�ƹ��CNrl���p��|���Z�PoN����b�:^����`|��y݋�D�Rs�_<�:o�����
����*D7��( � �����y�}���^:sk{��$������@���52)+ޮ/���v���M��d+H�I����6!�\�/A*�-2U�|Ś=��V�l�k����?4+�,�9���K�V�+�w+G���5���ep�]�#>06�j�9(:)Lz�1�! |e[�C�A	���e�"�;�u���Z�_�$�P��!�4�j&No���ۿ�(B:����X/��Ð���v��s����Ш�ej9�[�z��|������P��9Џ�y�����}
2N�1^Q�?��y��ѺqJ��s^º���<�ВpMϴ���%76��2��X�z�`T��$��l��>����oH*ד��e¶�i8v����nC#��׎P�AH��ɣ0f	���nA�SX��2�dLW�y��Ų�)yW�j>I���(H��ę�s�zn�٫*ޤ�r�@Q� n�;�������J�&	ݤ�;����I��AvA�&�%)3V�"$hyi��v�#��4�@E��G�>Dc�����b���e;� ���-1|z���/ �ac�o��e������	M�iֲ/�3/w����M��4P)~ob�����B%����nkh*_\�g���oK�7e�S�D�$�s�]Ǩm���//H.�\}&�Y�3f�-$��L�;�%,N�t�?F� ��D�;��X��$i2�܅I����N�i�E�(]����-��R�#��#yE�:��T;%�\�e�l<
�x����}�|�HhhD���*�14�"�Zt�.��"��7/�E�!a�L����b����qԅ*%����p��#��1P,>ӝX)���!!�DTn1��L�ra���s���[���M�:��v��6�-�^��q��t��V*�k���f&��W5Aʁ^QZk��̦��ߤ�9��0��mMr.p�L���{\��{����ѭǯ4�8[�)�kF��aG-���������qX럘��$ޜ�W,xǲ,,��pv�B%b�w��dȧ�6����$UF	0����\�m�5 (�ʃd��v8��v@'uj僬�B��l�,G�z���A��'D�.�� ��W���N��kR�t3^�l�Kv �=�`�0FuóNn�XßFB��B=@�w!*���m�p�B:�a�VW����27]Z�M�2Ӡ�%�-7����v�~�i��Մ}(t���AjL�,���,a�}S��l���𛪒�t����9ޑ��;��ϳa &&*G�c��oz���H%�I���dW� �ߘYޮ�S�Gr�����.���-<:w'J�!Mt�r�pf����[�<�EO���ng��Sy����ݩ_^��F`B�\���P��^�0�2ݱ��=c��<ם��H��a7�w����9��߫�����+����FsH�J�v���:ve�c��by:��}�7�!�Ԁ�gp@�v���٧�
:�p��taH��^~耭����]C��hLүY%�
�*�8$�Ɩ`C��5�lI�7�k���~R�ёa��U�����{��)�wٷ+E���;�
�lϜ�]�Z�p�
�*��1���u٫:���Wv��N�*4_F�(E��`s(/B� ?'s>c��lÈ�V���+{�:��w_��ZȤ�\mG	�|:����Q��H\�Ү�c;�*�a�4EFC��b�����~#��=T�4�	�b���--��)��o��fAa��4�R���,f���ٷ�^����Բ_��41g�b�6Qt&<3v(�=�c�k����
�������ί�7F-!y%;��]��A�s��e���fCy���jv��v��']aF;(��
��_f-��Y�P6F��~�pO��rH~�d��=�mnu�d������;�JX�S����u#�&��()bb�|���j4aF
j��ܩ���5Fij��ĩ����}�[WP�W`{���Q�pYt�d�H~C�u����m�`~��oCj@:7��]�ɻfuD �U���v�L�/��!_E�ۈ����/,Ӫ3����DnG����h����;�5@�ߤ�,怒j�XpaF4U|ɘ�3�v�n�;E��ZvM�{�.��v!��h�5l�k0J��U	T�>�%%�1�ذ�VN,�	��Ɠ�ć��sX�$B�fpx���i��y��n�j��w�����OJ_�W��^�&k�;O��9�-���`/ 3��c��n�^Dc�c��\�}����9�b�u�����@���"�ۆ������M�@/ԏ�;�ǆ�2yY|HX��N����R���EIW+��c�l�ki���I,�LC�Go�D�b��6��R�>�~c�F�<l';��8��&���LuOB����[�]�&.�������J"Vqx�a)�Frٷ	����A[����.��b�@1h4ê��:��0�x�Lf	����_L��>gw�B ����N�����LkzI�<���&�Y�s��
K		ߥ�Q/�8��
����܏\��f����2q�+�BhSa������eg�S0�@�Y�Q�+Xh7�!��+�3�K=�*ǻj��?�Q/e��d�Ί5@�W��&$YE��G#��_�H�J$EQ@�g�-��z�?PO���������P���x&��i�AO��a�n�d*���~�q��J�tk���(�-��,��i��.���8}��%��.%(aO{�).�W��� ��a��$ZX�"X��Q㾵&kSH⤺'��gە�$�!1]��ak����[�e�ګ�C����v*�V�C��JS=i�r@ϵ�c;%�����U3���ai�֥����PH-=��B�>�]s�i����<!���
��y�ɪ45�F��BƸ��$���5y ��ռ�]uv�o
^��jE�(���u�XfE �F��*�7�kn��c��a�<)�y|[����fxrM��η��r��Q�2�(�^�?&��=���7RX�ͯ��p�����z��jOߔ�c�6d:8����pJ{V	f7�OQ9�pg�6�a�ER�:�c�:���ҟK��l�@�������m���B�S�0d�h�B0�iqOkp^$��ْF������d�V��n���.j8Gb���f��Aސ`���h���X?�`���O��?�[\�q���,�Е��%����w ����
�Y��F1�����:�g�2��&{�ds"Ӹ������)�߳	�]o����`CY̚6ԙ��l������r��}�RJ~���G'�m�~�SOQ�_��'5�>�
޷�5���������;fC�g`MR�F:c\`��A�%���I���+���lq���l����H�c2�y>�AUw��Zjt�n��h#���Z�7"W\UJڄ|�8����;:�w�֙��Ԑ��)�V	�+7�ۚ�}�s.ktc���J���>'c4��w���Zj�+������,��5����o����Ku`�h�?�LU��.<��KR4	s �5:BO�E�����KP�B6�h�\�D�;o-�w�g����0�6E�+8%}��T�t�e�;�r�܈D��y��`��) ��4�w�r���xf���_��I�s�r_�nߵͿ@���B��`�T�NfSu��! �CN�Y8�C�v��KHKN�B!AW��ʹN_����y&T:Se2��n�K��g(߿-d�SJ�]�����6���I(�_q��7ؗNz]�����̐�l�$��3�!J@����o���nM[�)�:��ޛ�Ȩ*�Iv{��pvη�9�X��RAG���	%��\Í�f�e�4�؝r���c�;@[���@��z0�~�8����ٮ��U��*�>�4����	�zC��\��c���P�q��t��2�cI�A�w5l�5�r�Z"�Yi�z�яn���[�6��"�c|�qR_��j7q{�
d��Gx]@��������i;V����Æ���ߤ�ye�C�{��:�����m=pk���B[�/~Ԅ����		�yP��|�����;�`;�#\c�T���H�ԍV��� �lA#޵�ۗ��іoءz����d�o��r��f�ƽ]�U٣d����K�@wt/҅1󨪀�@�HJ�A*����A����tm/�t%�	h������n���|;c珁#y{]P�΁��Ï?2�	��m��[;�&�^�6�Fq��� ��M�В# ��;��xCj��F`��m���{zł���N|l�%8<�1P�U=���)(Tr0Cч�,�	;�F��qO����z���<�+�~����!�#���.3���Ù��sd[���,y����,%�	��,��Y:��)��p�Ku1�@JVW�J���4_��t����Kx�k�%�~Z��E$�P%��`��*�vy�^|&��ޖ1-#�/Xfd�nh�e���6��գ�t�� fVH$��{|�qP]���zN~�HW��t�A)GX:*�6�>}���1�Yz�k,N;�*˵���7~>��'��F�d8֑�h���e��N�@�{㫐�����Jl�-]wt���-Kx��T��Sʏ�ڏ�,�8�����E��.�H���6K��q���2}�^���t�v�����8�6�
N�<V�G��k�x�g��mm (ꐓ��������wV��%<�{�e�
�&uHƮ�g	�^� 3Hi-��å��X�1�/��XH�ynh�����V�;��Ӫd*Ǚ@`7�)S����z=#lt�G��6 X����zC�$>f�Xv����33�� W�>@@�Q�)}������>I��:N���n(@�T����btV$1xR�<�E���ku6��d7��I���F�UH�U�DӢ�jtk\��2bOOwA��=n�4]��@��3�[[�� �/K���I��I�M���Av��3[dE���%ʆ*�NLP���%c6��e�e!G�\@��1�Y (ŷ�{%�\�z��R�ok�sVQ��{'/s]!��Ӎ]������|]��@�S)�^��|SWl�h��BON�Y�6��eDF݁�[�ʳ�&S�wf��P�O�ܻ~�q���_0��5�X�<���b��o:�X�ԇ��^Pur�.Q���}Hk�>�N�F��RO�g> ��ܰ�w"�a���\K*����ӄ�/*d�Y�H�}�%�tM��zu;��o��X�R�75e<dlގ
/}CY�uQwu�b8���0�����Q @�j։� Vy�-�F� q�R܁���Ƿx�kԿK�j��n�&��)Y�G(��+4�{��#������k �D,��f����iq����	ꑵ-�P��zPP�`.�-���G|���:Ǧ�8��UTS�I���D�O�ĉAhlq52`H���i���NԈ�Q;hz��G�Vl���"ȹ4��#Y��f>nJIL�Ϝ2�L��븩��)���/{KᎿ7���	�q.��k �i0&A{�{��q�LI�6�o����+ce!�Q����&���
��ģhCa�昵��c��T�9��FQD��mC,M�������1�-qA��-AF]r ���	�����X�F̽���[r
��ޙwW���N�6�D����w����G�$�l1n�+�d���|OTyFN�� d0sN�t�7�7GM�%Rf>�g�9�kK�a&�e�?z]��J��Ĕ�.��߄��Z�a'Bk�	{
�*J^)��1��Ɛ9��x��� ��p&������x��"���E����2)�	Q��� @.��2��4�m��j��G�eC�L�3�-	u%<�)�z!�#�w�_fU���4䊢��ml{�����Id ]�����.�$��#y?\T��z[�R�tTA���tб�pJ����?�s�[��u����9�t.�Ph�3Ӑ(����WvS�:A���j�l�Yl��`�ѭ���F���BV�g�x2;�=`���+$e���i.J��D,��7�Gy��`@¨�-��?��z���5&@��\��aUF6W@����*�=C0m��~ǡ�㶸B�⩔.�e���L^�\�RW�ػ{�P�q�]&�č����w��f{�{�w�$��ܿ�g�zu�(4%N���(a��<�:Ꮹ�/9�\�RW �O R��*۴;����� �FYT���	�K�5�U7�,b߮E��遲��7;�w{�<t��!.�ZS��rK
�ʄS`y��x8�2���3�ň�����#���8-�e�V�ZI6�2N+��'Œ�0�C��+Q���1:7�.�I.wR�U�)鷒�'�}Bu��'<���(�Б=* ��e��H���Vڔ����C���uS<�V�5H�
��r��P��Q��0k�����K�<T�(�'��~�
uT�u�t���J]�C���sŇ��2�<�.�G<���1(�6 ��G,ú�IW��e���tz����^i�4�0����G�B�Op����r�e��܊��7�재s��{�=� ���[sM�XӾ��&y@��v ����5�!�Vx�V��b\Al��{��7�ʱ�7��8�·���[4�9ہ��`��:��D��q����`�����WIVh��F�?��c���������ǒ���T�J���VhH.������5x��Y�e�~!:]<�rtyQld���:ch��w����;ݵ���u�o��8�h�@�oV�vr��;���B:i��i���\�������/X����KY�RAv+����M�5���Wx��t�y􅯰r� �5��82�+1I~� w䣝0��*�[w|�Za�=Tm���b&�%�[�B���)���;:�ê�D��߅�	�.	�\]T��m�>���m��"�ݔ��f�S�&�'��H,6�� �P�]枞��Q�����8�`u���UG��Z�Y��0�fl���>����}���y����TUV���}�Z����3�I��R<�a��$��,�T�BG��=��Pɽ�^�7oK,�o �:�,;k�,G4��d���E��_��c3�lh�"�B?�أ �Y�`�8TC��Z��{ )���k���:tҳ�db:��=F<-v��l@�@�Z�PW�v���[m@�E�����!�K1�Pt�%pq��:D�}��z��z;����ՄW����؇���p���[�"BD��"�p�7���J��;�''FS�����?9]
��=�g�GQa��<z���+��Eb�u�����R��٢C����������v���b�[^j&�,s�뺥�Z���I«+0�Ad�h�>�aFK9�*i����њ��J�濟,M�W�|yޮ�����8uw;���y52�Vb.�1G���pA�����DT������X&�5�L��+[�C��i'3h �k��1�{�#2KЊm���L�Ԗ�=D8����y5��O�-�g�6�k[}l|�}�,�{���=�E�Ǣ�YO3M�Hp��T��͠i���j|y�^����?��u�E2�����c�<!�����m;�*op���������P&R)�7	���#�q���$ ���{$�Y� 2>!��ê�(����2E�7�b2��_��gkr�Ӭ �t���<�_�2�K���Y��Z���$�������Z�;�	(�������h��2.�|�SW8�:������Q�����tX'�F6`�#Q���Hy����3R���a��<B!oC�}�/�x5����X�7�퍕�$#+;���t��Q����! ��Ӓ�J?�-a�"eƆ�wct&s�NV�ȼ.�G�b��@�q;g%|��J��{�D`$�c��}�V�n�k![Ώd6�Ξy[	��J���!��-��Yɸ��b��!�D��!$Z��t���S����9� Ʋ�/)?�Z�!��?�c*���������b�A]��;w�A��av�WF&tˉ���,]�g�s���_�u������lhN��U^�u޻:�rk��bX;�XA��/���2D�����]�p��sp���$��$�& �u�la��>X�jH�{�,��������~�oW�`�N���ף-w+���绌mZ|
V�p���4i	�6�0Gv�22�I��b���� ?M���-'�VhK��XL;��Ԣ��9�8	�Ousv��SL=,!ނ�d�.�q#�{��V�@�����r/�T$٩3���Gh�m�SoR.f��Ѣ�k#�1?G����<��H���INe/t57��N3Q$f������+�>��y�C;e*��fqԗJX�*����{Iﭸ���5)��`�2���B�x���D�Q�4Ɏ'֙T �Ͷ�d�
�#<7� ��b�������mĶ �'������@�&P���|�`F��,��+Tf5��1}��2G��Ϳ�4�x�����R-�$vm|�[0
D}e��d�o�	M��%G��O�Ƴ�Q���3��'7���C8�9�20�Ϲ<υ����bBx<�?ݤ�4Oiq,��k��03���6oIP�4�Z�(!��6�7H�L�w���0�~ʄ90=��o@�i�pd���2��&}��^5�k�	!��"Ď��T���Xr��r�4�-j���
�v�������hH�p�1p��K�E�X?ɯN��mVܬ4a�_��CςH9�UdI~�\�G_�Q�l1��b���Ѧō�i���6 j����;Ͳ�S+�}�B*0�}�h�ُ0���.n`�$�l���D�F��gT\M2~=Ƞ�3�u���:���lH�=�A�1ޢܷ�/��tM��L��X��ޢYV��H]�)��� 7̏.p���4
�y���^(yuMD�|����������M����ug�C�����O�"��5L�o5Ôd��Vtw�V�) Ƨ�^c�'�bD1u�:�G�̠��uR��󁹇�;img?�Q��k�^��9��Pl�y��K��z�0vr�H�v�p f�$�^n����naY�s8ҁ�i�(l�%c���E� �ЗG��ZV�ѿ@4�7ԗv���U�a{Z$V��h=��l�(�R��l~�+Gᐙ��`�6Z�Gf����M[n�nyq��e�����Űs�Zԛ�k5������m�3\{�����B�#����G}�����:�{2kz�Ⱥ��@�����g�-m�k��?��
bG>��ƈrÇrU���	HMJ�5�?���l0��ɨT��q�o�A����:��B���j����n����U��S]熏*�Meå�����4����1��8�h�H����zpu�Jt1#w>���$^C�y���EcаH#�s/�����Es/^���_v���7{������sS�OJaUZ|����;=�9��P��{��bM<��'"h��1��I��hR��s��5�vG����~5��\�U/J��O��2- �V�Gޝ�oY؄t����-���gN����!���Q�܀�1�Q$� ��HX�<��)S7���T�0��r����!o����3[^��u�vhc�65D�ܡN���p��� 7�RB�O��r�y�'�ʜ�y�}?'�o\��h������<�~7!���)�sf��Sy��? 4\'�����
x�����k`y�h��C����
A6�;�X*�ػrs:��!�$� X���fɡ&ґ�SS���#DL}�i�8���`B�@�+�w��B�UԖOĸ�6�b14Q��.cl�uH�����.�3�(ͽ �0f-8$�J�kr&�x�>Z8`����x�>��':.kt5&�����v�/.5��ڪ�4��9��ߟg=N iRe�yze�"mm��B���m����� ���ȾV�> �!�\�P�>Ɇ��4�s%�U���� ����	INN�ǊyU�]�f�1��'�����8���P��Ig��jn��q�	���n
�����|�*iy'����/OF&���T�ɘ�ձ�e� mb�ID�X�����y��$����C�U8�)���<ij�!r\�$^�n�&F�r�R�`�-��'��V���p��0��۾r��0 �j�}���й|g�9.½���?�@t�rRתE�>�g�p���Y���Y��ʶ�Q��v���Iw"�M���GH��mӓ���KB���d�ל#�<��}��d\o���f}��_\����Z���xaz���n��/�~�s��{��#��}�9��)L�)"�B;����S��_*el���V�8�J�&�	}��L/�E�A{<>PA�$���}���1E\֚�v���R
j�À
_�����1ہ{z����G$T�'�����P"�����ǉ��e�Bs�!ɥ��]�|F����`j����$�m9�9�\�kY�n8� ��礅����K����O~��pw����8$4�˘�ɜv��Ўw����m��ck�-�ϊ�}ނ:u��v���U'`�z9އn��_7��c�d�V��U����r�bOo�$-jy��܏��6�[��iޥ��q���vޡ�v@��خd�OI���G��q��K��7��� 
p�?��iu�8��x�/�/{� ��q���
T�mq�T0���e;WJV#~S/���
�Fx�]c}�f&ٓ��h��t��vAѴ��!)�[�[�
R�rS]�ߦ�6HT�yIo|�9Ә�8��<��A�r����r-����T�6"�fѓ?b[��N�3u�ir�<��PZɤQҌ��*�xv����*0�$s��<�e�D�QZމ��;F~6��ۛ��7K�6<�c0y��O�6���/�(.�;��zĘp9 �^��6;�T��j������U��\pŖC!vؗ�PFܱ�Y�}YB�7۝].�[�o6�5�dH�|s�2N���wc�"���/K1�5N�l\ �����Be`vYA��A_Ѫ�����w��\:i�uVl�/'$Q���d=#2�d�
��bZU+�oyվ���n��7_����;m��J ������b/'(����<p�:�Υ4�B�q��\^�	J�k@��_�1�y���@�)2��*�n�^�m�ᘙ���y��;�Xt�͆�(�N���#��읝��Ő���ɐ��i�n�
�������=�y`�VݟVi�+���چ�(��R�=f�@�Y��Pw1%Cq��-�����P���#�&��D|Ss�@�yk|��-P1\�JZ��b��[4>!�1Ӹ�rQ�����@���5V$�Z�7��{�}���U��K�*)Ob�+�!^L�~1��r��81�#��#a5��9�J3
j���j(�K߽e��7j�S���f��ꃁ�� 
���\���΀�ц89]p������NX���:�(K��EC!���u��������#FZ�"�δ��/z���wp`T�ϊL�/�� ��F:S8�a&�E[�x��m!�ZisP��4�:C?y^���;��1N��埵���9��G�VB+~��b =9�t޹�YB~�zfӐ���=���?�G��\���p'ǧ�o���ߪ��xƷ:)c�p�w��J9�� /1<�,��������s���
���B/@@��hkǋ��[���P@K{�)�%�m��w��ō�\Q��kضx�$��0f�M����XGj���D$��[�#���9��`�{$�>82��V�������bf�r3�\M^(\h/y���h�
�Zܴ�x��E|�����ь��`��]���sQ�	�2�I1<ﺪ'��>�|Pb�6m��c�ر�.��䢵aTw߄+�{yó5g�_$C �.�������Kʐ�{!M�@�>]q�m�CΓ+����Ʃ�;S��M�q��p��)�|W�E��[Gef�K��?6'D˳$w���(o���4[��nv���E���z7�mT������w��K�2訲�g���0o���mZc���k1���Ygcx+}t�b��r�s�X�)���2s^�����ߗ��0�H~�8��o%���z�i٩���}6g�� oyn��w�i�N�1����n�AU�ƶ�Z� KY�`������W��ړ��#\�0���q�>���j;�"6��3fޖW`�����}�p�M]HVx��q�.��֌2:��2���q΃Pj9� ���L��3���L��U�wNk���J�2��`4[��T�e.2atOSjb���l��ޥ_��GO���o����S���-/�Ή�c��.�4�ݤ���A%��[v�"ݐ
���~��@8O���E��W��6�I����gmGx��a��Փ�Jf<59�	�E��J��}���qXN&�j#�S;��*y*�JP�����Ǽ��c��T��_ی�2r�������gi.��Y�3[`��|� d�с%o�nV�*䰏�_)nKGĝ�g��c�F��4!�_|�7V��~f����'�ު�YP�ڹZ�Q���R�ȸ�>���]��8LՊ`��s,��Kff��a��Lv�&�_�4��ڤ�e &w���Y��woD�:�gxnY+��W�fb�e�H�>T;�Y��6��
w({Ɯ��mi�����C^f��A(�~o�;�7������',͒�2U��dB���3<�v�0��yЋ?h�����Ww=��c�ڡ��\A�け�6Θ?��c��?��1e(�B�ULf��%���+S�f���`�
��c�ŝR�w�'��e��މ���S�9��@�]J���xԞ�2�����
�0���2��d��d�L׈s�J�<�-�h���R�l�4��Z��e�)Θ�\hϕ d����W5���;�Z��o�l^��P����-
�'�~��O������)�O��o��Gkr�[m�p���VKa֭ 3EʹC����)��$>m����]/#�����6�|_ �ys�y�ͱXz�5fSag�$��p�8\�J7'��"�E~#��c�T�^����b��Oq�y�;�-�_���4�Qܡ�Q�R8����qz"}U_J���3ZB����ְ�w�lc������+�����2��f�ul�Y�-L\���>�������
v�&'=��+C��<�WHB�>ݙ��8�b@�e�@�ly�gY��Z!�.m����j��̱��_��&�P#�X���/J�0���%$O�_�P��!���h.�S��J�=͙�"���7�@j?�9�_���\E@�b�?�1�]�a�X@_��������$I
����ؒ_�1�R�߷������\$*C�x�<WEٟ��j��_��\������/06d2O>�Lkp'.�'z�W���Y����%��Z�Ц�T����.���Xu��<��wt��"a�}�I�/�E����Es�'���|�"_�����`��&*{Ĩ�B�:����&�) �U\:�*����0��a	iBI��^�D3� i�>Z8o>���_Gf���[~N��g.�D��W�j�Z�\�V_��"���6fN���3�
�*��Æ!$�����.;­�~�/R�$�M>3ǻ�u�r� �Z41n����x'�˻�$����W��&�&�^ ;���05Yy��R�x��7��}P��pP�/�%�����3PM�#���gKU"gٍ��[㨂:"���z=i��lJA��;�ou��)�8F��i��$��JhuB�c�����[K�4@1r�cv��'���_�����ބ3��$Z�j3����=��=7.Z���ww���u ��J���b�_?[-E�8jv��n�m�̡oj�<i��#�i&�g�c�ۥ��2=�I��|�iѽ7tx_!*��S ��e^e���!��Z+�_`�go}�"��j����{:�@%M���dgQ$�WXם����`B��	�i�a��F�U���`����&u!�iQ�^̺�_C�_��Ǫ�o{"���2�]�д9����Z*,4P��7�}��&����.�~�q��}����kh� �(K���cm�>7<�+��K_xa�	'�J$-	����Uu�ӄ�=%�'�gg';��t\��f�.ih؀:��fC�;�yd�/�3r�a�4����K[!�<1����K�i�F�՛�N�A"]�
��o���7~��n�� y�*�!�7h�Xo�y1��t��2�@V�>�،��_�`z�$'�0���*Ә"_�0��Ofdm��:���zH���2����v�3<�Ш Dځ�$͔Y&zU�1J𤸝W�Z�P������C5b
�mUzc)&P10æ�-�P2|؍z ƭ~[�3[��b�'Lnj�yC��F�����}�/4��E���|݃"��x�b�)״Z"�����p��c�Nh�S��7L�S����2c	-&$ȶ��̷����ް��d���goi���455�������}[EP4��m+��@�#��	�N�Ƚ͋��~��':�` ��)�~-kd�¤9X�Ô�r}6*-�qw��v��<����J��o�蚛>�7+ �N�V4\���!��A��1��ߝ�Jz]����)�J��W��1c:����m,��>cŝ�m�H9�TI��ޅx�����>I/ް^�%+��u�i;�ےxȒ�Z�z}U��*���&�)��N����F�H	0^ԱjbF<9(����gy�߹���||��ٷ	o���(�>HD܈6�_<�9��z��x�Hgp��]���(i�$9O���bg�ٱO��.k����x��q�f�"lU�A; v ��}X�B�N��3�e'�D���+Z��:�~B�%��fL`����̉2��vl�
X�B�F�PG���9�	՛N�\q�FO4�a��0����\�m�i�n�<8�Ã#����3
	�֏"��ۊC��ވA�ҽ�p��&��N	�n ����zHT���s�l�I@���%h�7�%�W� ?��I��(�xK�A(�ehs�Z�����V����o�d�ű{��9���-��.̱C�6� �¬���#E9>1/����ׄ�5�Qw���#��=�}��׿}���r跲mْ��&��^�z6�����z�!�a#�͙�t�+�
>�
e/ş̂s�F�G
��i�l�@P
]��w�4�bqR�JH7I2v�Z�ħlܜ��y�քKm�.�����Q[#\7���V���5K�f�k6A��
2�d6?p��<� B�^��+"U��
����LJ�'M�in`����s���QZ�i����$���89�նm�NJ�1#�	Ƃ�.J��]�l���WqA��ǃ��\�q3k8������e��{����eP�I��.K��uu���^�
�qyQi�Z��}C!lٕ���.y��p�T�8�鈚u۳���%��*t �rݚP<����B��q��=+͍|�����c���<7y�1�t�d8����E��˔W��ƻ�4����rg{�i�gP��#�Q��
����w�9Ḿ҆\�i����
/�Ə���g�xh N)�&��.���P-��P������
���p�
IE'ƱM�Q�C���#��2����
��_U�D�^�q��Q���I� &���xl��8��ݵ,MJ��*�yQy��Q{U�l#N�"�{�W���B;e5���]��kG_$6O\Vu,�H!�4ޤ(k�����b�{�.��H[�\}3�o�`zQ(1�4��(����NE�y ;�����Ü��M���%�Oxq]�$����X ƀ|1�7,�{X�Vŗ�Zj����(��)j�s��(��6��V�`�ܡt�3��͈��G�J?>6#xI����tQ�ܷ�]r�q���	�rJ�7jf��e�.�k�:�Fq$��Y�ڤ��Y��IT���jC^��r&���6b�a�P�2cC��ۂ���ْ��]|*�wX�; ;Og�L��g�ʱ�ZKj���k�Ԧ��6����<W���p��8 y +)w�������kK�M�4�EW���5�7��@�Co)��6&s��<�*�h�E� �J�l����Y�[E��D��L&[��,��*)wڅ�%�!J�+%��޲&���T�6���L��E�@�r'���J��.m#e��<�H���@[i؜��S�X����jmlIΘ��2�}}����,���~,�k���­�[�Gu�-P�N�3���GX
t�;7s��c�#�@+�F%oJZI���xG���l#MAP6��jW�̇�X�j���ʐ���Ev�"��G_"��t��,vK�y�x��M�;�'�.��R���	����Ȑ�w61C�X}���N\�;�$9�Ը��:��E���qV�8��q��q�1��8t�����
�}J\�;n?�����Ȁ�6��O�	Sh��
��8nz�ُ��z�ա2����DA�j��&J�b��w��k������1N��Px��	]��0�PJZ_��˪�&��+P`�>=�{B��N4[�I�(_�a�Q�uS{&��q�A˱�W�[1���L��Qj�����ϭ�x��Uo��C_�CJ�I���r��qܒ���wRm2; ��5�`'�"b%1<��ٯ�`�\4BE��@/ػ�8���-�����
z�Or��n.�/�y�m�k������UzU��Do7�ѡ��r2�F�d���TEyM�S*/p������n�K�!>����q�m<�� ��U�Bb�}㗭�l�(�����.�(ۭ�̂o�l9�ҳ�d^&���`��BB1���bGG�r�r�,�d�4�A�b@ �,vo���<�-�?�I�� �$T����ʡ��p�	�=9�C���p�B���M�e�-�':�
h�f�¬�U�(��yLO:6\W�tW%��������f��>~|��c��N�f���D�_�kQ���t��k0�&��5< 1�`�4���4Eyez��L�T���Ge��D٪W�5�cG?��]�1�m�R�g3R�P��(��)�Y��pub֣�5�-�����Y����U������ѧ��/��,o#���k�)��ޓX�E[l��hc�d9WӋ��m[>٨+�ĳ���<���|k�#�(�����)��$�"#�z׸3�Я���=X\�c��y�i+.%�1,��}D�H�"M�(���$�L��nKJ?;��ǟ`�F|E�h��U�v�/�౵��/���䧰i�~>����C�Pc�H��D�)\2����Os����4�A.?������1�rҧܬ�[�K
�hU(��'��F��C��C�l�gW�u8yG �耂<�,vP�sІ�7�v�\��*\�@ޟ����Y�'�48�4v4޸]����aK�ׅ�zܐ���V���e��)�\���=�(�c��M��w
|XCJ��2?�=w�/�<�_�o��^�7��"�); R�?�zg;,��|3�*��]�;i��=)�,�؎^~)�����dT������i$��z	^����^���eM�.������ЛA��x֋�&ښ�\�(��&�@W}�R���0NrS��}ۃ�Ei97��z��,����������C�jF���h��9��}��p��O0�����:�$ةU�\Å&�$}�8�:w]�L��R,���Y6�.F�e���s��;�m�,e�\�g� ��?R8���6�״'8;�S�%5*��~-˔	����!�Ső 'Z��i�{+������k�2-��i:�wD��nE3�\~@<(8����Q�����ج<��k�����P�֏��"u!p�'�l����(G�ޜMb2ǝޒl =*�oI�=��|�|zT��(==P7��S��� ���+r���6��&YiD�U��AD��<8�L!���buy�L[�|zd����-�ݡ9�V�JK�m�RDG��o������=`��6y��\��Q����TJKd�*��-&3��A�y�fc���.h��;G44ݐg������5p�<�5(�]tqպ~Q ���h�%|,����{f��<�1 M�+ox�6�D5�m�]�l=q���]͡BB�Nqy�|*�nh�o����e!��ہ���Y��Q\:�B���J�Rk�f}��������a���E���n���%N���G�ci�g+}��E���0B�C�x���,m�Qz����sG�x"f��p�z����ۄ�+2#�����g��VF �߁�Qw��mj�א��.K\}T�K����`.��Q�Ym�^��:;�MR�Sc���d��Meu]
 ���\��m��Р��� �q�e���%}�Cl���%�����Y�7�Wi�`����j�:V�W�����-�fM�
b=X��z�#Ӻ;-m�"���E���p�W�������%`��>��dׯ��jH�+SG�-A�t�{��&�@���B#]x ׹���l+@�~�{h�n�O�0,�km�3M��K��*)��5�/@���O������!��d~�"�͆I��������#N�j0�,)��)A=<"&���"���[-ӫ㠞=��ךּ�P�Ok���bk�UE�����"vjxЃ���'%��s���Ro�l��!].���,�䎞i��{�s��]1��q�Ǝ�`�3_��i�j��q>;�QYE*����^�LX�;ԅ�����K\4�R�v�Cp��e;|��ފ�c3ƶm�`D�>�ۑOCxU51g53�TW9ޠ�X p��<�*.�]�~�~?'�_o���<���E	ӟ)98��ŵn�t��Y�i��w�Ԟ��E�ҿ��ļg|�@��CO9s� �o���
��(/�<���zqmm�[-�f��o�G�t�&�P�$��b�s��:���O�����.<y�H ��z�3�>2�<�,����c!,�Є>HY��
J��c[���r�kP������+%-*�|'3قTϯ��C�f>�C6]���n�`ǣ5������}��#5�!��%�,b���V�0+���`*��[v��B[�Θg�^8E7{���&�!Ǹ��~� ��߉��,�4<Bx�"����5�˥·���	��2��x��V��=t�S/����`���\�!L��r��>���0��{�O��Rcy焠�ךq-�5W� �� s����nxH�.~II.3��-Z%5��PPBYO`p*���t����$�]
��
oy5��_k�o8D�x�����Z���]c�!+�ݬQlwKƞ�X�x~�w!�U���qf8�O�ǉ��wZ+�-T���g:F*"1���b��N'������'��&w �z,?�]t����40K ��H�,d�-nθ���e-5�����lo�:��.QT�ޖ귟>��v\����j�_?p��˽5	Suo�~Վ�R#��A�R�"�r���w��<NvY��X��:��#׻�_��c��:��P��$���[���X�&�2��p�q�{[�C/��,�>��l�υ�N2����� k�ys��3U�QO��Xf%��=k��ż�[�t���ù�I�e�yJ�r��`��G����H}��ּbz�����L,c�tΥaf����aFpd��Ou�R�����Eސ��̺�o�/���Z7!b�Ƶ�L��Xu$�Q\���C��Ɩ��K��C�y�.�?V�
֦I�̸��/'0Z��ʓt[�@�����C;�)���4'ug���2�yaH�,a�R1]b
���S~k��3����k�0D9���@\�2y2��d%��,��C��J��~�y.�a���LU����۾����������|���7H� w�#��Ȏ"75tG�S̿:k�䳉�v���E��t�}��/�� ��]�=v�t�bэV�qͱ�t�E�H}�Y���WPq��Xﾉ��T���= /�GA#���C�v�R�j5�[��M9��Nd2
ѿ�2��}�"��{�M�;����/U���S��<�:�89��4�8+pV/��(�q'ⷙL�lY��am�������������*�g��$�MCuk����P�@_�VS�
��|I�J�XȢ=�z���>�r���q�8�p2��(�Pڠ���'���!�M������	{e��nZ1xm��� �5$��1(����5����ė2��;c�.��Wģy14.�L�����{�T�S��є3sǛ�/��
#��F����)D0ΜZ*Q�� Ƽf��^��Prg.���v��8�i�����_�H�Mf��"�f}}�~�*g�zA���}��Æ7\���I��1�.��>�P�k�9>���I�+��?�	�Y�I!o�Q���}�����q0͂Aͱ�wAxs	
���Ղ��0N��=�#�[���iDn���4n�~9>�E�JK7ߊ��:�`�V6��O�A,��z���i>���~^oH��&iw���q$����g�U�D&����e����7��D!�i<�yE���U ��Hԗ��De�;�g�����%t�A����eq��sjYY�z^h,p)��8�f��CD�c��<�̉��?�܌����ir�V�qRn>��
��lq�#�V����?�VI�����r`��*��:uȦ�x����5`={���UZ["�Q����˺�zD��|��n����V�i���N3��U..Ԧ�_���PF�c�^�Ώ<+��L�ųQ4��Q����N�A��qGg�og�❨��\�Xn�gZ;�n@���GKP{��7T| ��c��J�FN��ojD�o�?��L���'DF
�6w�9�?���c��"��=��.��m��,���}�A 9�å�Y������o�{EOq;���U� >r�~I���K��?(���cQdk� ì�ܟ�kqW�����::������ ��@�cQ�>@V����l������w�y��b�孩{Hi�OM#�Ń���\21)��9�A�+:�<o�K���oK0>��\8w�"�h�� �>�A(��+
�9�~�~a��_���2"hνu���:5W(N��-�oݒ���%W�`U�=٥E���G"�/H\��[�n˧0{C�ڱXy+��46haǐdIzQy喒�8��b�␠����`�jg1wc���9CK ��c?���S$	��Ѩ&����P�����v�����H@��	�h�a��t� ȣ7@�}D�~������7.�1.H���)���&h��,�5Z�����00�?􍳔��9�]HN=���"���F�ɺ��0 C��u&�GYR���^�Q�n@��o+�p�f2D�RP� �+jNd�������
��>�c��Zz��%��k�4�`�A�z�E+)�(cP?=��ZI�s���9hMɎa��A��	9�ΘrH�TϪ��a�� ퟗ�4S����b��|�&��!��y���DuI%����/��eް�4�I$�<�u���5�;\����	m%i���|q��%�P�x����49����[�6����"��y����r�c(��^}O:�`~���x�yU>�ܐS�E%�wr�nx{q�0�ÛnVO8���&Vۑ��Ҧl�)OG~�n;X���[S�ũ�*�9���ǎ �����h d����vr�݁����FH��6@���>8�Ƃ�k�;9�z���c����Mu�a:�6����eU��_�����ս�E�I�ʸ����ΥY�F�h�P���� �O�Σ��2�����an�t���Oݙ�U�#I�HS�$�+��o-��cM�h-Y��XME���G	􎈯��I���b�E����ycʾ�=AQ��V�Ax�ۄ 5_#��f���̇�$>C�.�!if7#δ��!_i�_�v7N�q���+�M�.����W�K��U�/�f��W�ؾ���A���t��+o�\E��W�Ws@R����_nu��1�Yé��g/��W6�����"�_��K^ŧ��D�1S��\��u�Ďm�l7���$���i&R]��8a����{�\=���R�{W�-.�����\/K�f����Z��N&�P�4�[i�vP�1���������ڭ|��V��] �g仍/a�|����ꢕr��.��L�D	O�����GEf��l��\�ۂ��M��)�4ۑH�,��`��;JwU�!սIO�__}�_�v��}����)���}0��[��֚)��]js�<�>/䙕�ILY�@��=�e�i�����|bW����#�7��G���!�Qg����hE�������԰�<��Վ����=�}O��ΰ�;k!�	��Ev�#=@�$he���.�J8��_n���X&�K���j�J��c�Ew�`�7�Bo��7�P�<��3-�|��])�)�ZǺ\>�C���a�?����h"6'$���:�:VIr�m��Ca8Ȳ3�-����z���ӈ(=!PF4@�"���;�Φ�ZHDV5a*���g
�:��o�9�Q�B>#ޯX�2�.q��~h~�8��H��M��Z��ֈa���sb�ʩ(�k��a���2hYf3x��׆��vݨU���?�`Ȉ��9ݹ��$����s��,�ְ:�Q����*C6�J�aLh����`��=З9����(��o��!���&�[��|l&Ol�=�p�џa���kpV��ɃL�7a!J�����߹	�T��̆�3�Ndh�R��G�KI7��T�k�rk�r�p*,�s��u���q�D�;��)ˋ�ܖ��iJ?\�Ɲ��J���21�(&O'���C�K�V=���QT[FK��_������rۜ�!�"�(�c%�a4v�~��*���_G^�v�����b��d(�q?]
���Z
+*�RJ��<?������M >�c▸[��Q��QDP�H��9�t���)�G��l�+\(�~�������$��,=��]t�/����͞nDIt��]�W�����J^���'�e6z������_ �d���n'E/��r���e�Bw�N�k4�������d�h`&F屑6�z���o:	b,St��b�j,
�@�8���7c�R0D���k[N!�z��=�}���Jd*3��[6����� l<~-�NX�p�bj�5u�|�(�K�L�˄�o�t�q�-<7φ��j�^�>���>��6����-}L����������HYO�/�PY���{�i7��[���=|qva�Qe�G$[�Fh[���|�$d�
)��Ҡ�e_����0N��8���(�����0((��d�g"�����-�M5�3�V���)�1���=�$uHܹ��"�GJH]I��;�dď�Qv�Q���4��C=>W��ux-|�%�$cB]
N6��
j�4�����Y޼hO�[�A-
%T�(_���"�f�m��&��&#o�vGyT����~e�0
�]��&�4�����}9���W�5
߲E��	�fl���07A\YMVp�x�� 8���BPu.���h��Ojpڡ_%4V/ak�ڙ�[��p�����|�/!�W]'S���b�N�D���hI�O�/gM2f��]r4�$�q����[��9�r �pk^6rs�WJ��|���Z�42�ф2�ص�)-�	�Q��N��(��ي����(Hi�#!��";�")�����Y������zǜ��n�4��|�ว�.��J�N³v�B�-X*-B8�yK��,�{/ե�b�[Oѡ�l�j�.V��"�!b`��M~��������>o���X�;�����>sR[�e��@ī����_pB�V���rG)Q�+�d��x��o[	:�72*�V]�Z�{��9кvU����^���z�Lƪ�o%�Al���I��~-�e�k1^ېx��&�V�Pl�*-�W�	�#���Zb��@Ԝ:ƶ��-/�-_��u���6���ĳ�e	����:���6�q	A�|w�rsi5F�1� !�����茙ݛ���4mS���%�kQ�c僉��wj�*i�ת��!@(iH�ڠ��4�>�?HDT��J�F�-�F\E&��^����s�F*���dt��.�ec֧��)2�F�ߙK[��CQ.Za����<c)@�RpS�;�p�1�}���I6Էa$&�/ HUt�]���=�^JDc�	|��k2���y���C�-��!Ϊ��Nر�θ�����v����8�su��[� z�r+
BpOQr�S+��m?���~B����rE!�{s��V� �Ln����K�-@a�Ԥ]pBC#+9j�� ��egriKG.��*��j���O^L�!b�	���6���Y�Ӊ�V�x5ʺ0�b$�C`{.�\=�'Q�� :�^Aݻ�=z�
Kq�D����3��0E\�ȏNS9���|H�K��5�����5�D��Ng�_'����#+=�/�!˪�D�8�8��סs��z;�V�����.�B�3R�3sNI�酮�&�.WS�Ų!W���{�"h17B�4�j$��M���Ç�Vug��be���r�a�-X=�\d�\�Ђ�.D�d�,��Sgl�mE�e:]�N��D�tͰ��v)���ʆc�v��_(��b���6|eӜ:�%�]h /��YH�8&F3;���IB��:��3�ih$d�U�KIk��*��Ҡ"VZ�����,���))H��kl�B�7Ŭ8L탵uȡ�v���Q��;�,��~$ ��IV=Z�RͶJ
<	���V�HDK֊,*��}���۶�'{���0X�TN?��wvcN���~8�ds�^k���	��)/�rve�{Ox�cg���S����@�����T�Ћ�X���ҝ;`Ty�U�+��e�X��(�@��6p�A�F���|0�ߢ���0���t�DS�r��a�&�"=�;�Iڴ_.�@�%��A��3���e�R �
ع��mW�I�=fN-���E����2`��h�F?�'jj�I�[��ֵ"71��}�����;�fP������/��ķEI���GsQ���gzR;~هˠ���D�ﰢ쥀�`
R�W�{�g胚�����LV�&T%q�j�"�8]z$Z��cze)ї,~�⼱� H&��g��ˣ�����-K�<��y�br������?n�F���"���� � w����JN~��׺��"sW1}������#h�Kw��V4��;|�T��P-�W^=�ٶ�b���Y46���?g6R�PV�يԯ�o�\��+g$l�'=�ఇ����r�D�6�av��z=�,�f�z���89�/��6�D�v��2�E.
يI����DÝAT&:�_���pEM&XHg�(s��p`U9s�S��
��[�&�/Nz�C/`Y��;���
im&à�p�2�U6�D��ՑV�3č�
[?K�R�A9�#$�1no|	[w ��M�� \ߨ謔R方'q���.�k ����
��k��P	�� t�X����$a�y���^������� Lo� [�Ie�O�Ĵh�^T��m��'~��:�������{p�Gc)�5����X���,���"0rA���H|��ٝx������A��A�_�|㵽J�x�+�'	�m�½?�*��\5��61�n�691gj�0Mm�
��g�NdL�V�Bs�/(�[tf�bE\*xǊ���ώ������TXU�.�Л��k�3gF�Q�~Ǒ�4��@ d�BX�_P�9~� ����g�P�!�.�����B[�'?7mV�D�������Hp�|�����h�%�E��D���ґ�5-�;:r���f�*���f���N3�L�4G ��T5�����#"CHv��xJo�"*�lZ#|����,u����f�fN��Q~�	�G�|VxG햝\U�[b�$����W�7ul�Q�]��U*Gkm{W# L����n�?��_ƣ0�n���DI���뿁���U�s��	�{��-"U�&��'T7�-��I�{$-�m�!c�gg��RV�'i7�<S�<5����@|p�"�QWe9�ĝl�R[6;���-Q%#J��:⍮����+�=����6�.F���g��@�߳��F'��6�[���Y��7xF" �?է�N�|lC�u�7���T�l���Q��p�M���=ׯ��3��NS��F�Ԭ}�j�vp��$���o�z�&0�E����#��:W��1ę po� �Z���|P�}b�$2�|�Q��`�p�&�k����2f��xC/Z�ߗG���"�Q�?S�h���n����@C���iѹ9�B���^��
x|�-�����w6]Nę�<�~g81��1��nB�ROxk�cp���ޚ�ݧ@
��o�"o�H2T	
�w>��@vr�j����y�I�W�z��/�����%��v�6p��,6���_����9�ikD���r0x������g�an�ȗ|����v���vE�M�h��DV�ueh(���(�m(�ֱ"�nk56�����u��=k�UÿJ�x�2�-���W���ȣ���h��{�f�.����ж�p	�����Þs���p=�c�A�\���Ʋ��Ҹ�a�k@ô_�o�-��$��tѶQ+Ǫ��	0� Up˸������n�7L�>n�4Z�&��9M���DU�w#`�x5��u��Mu��OV�kS8�#@5 �)��|69ׄFىl�n�'�+�c��Ң�gT;g]��iG`�1e~�w������<9���_��\�7�*,�
��_=>�l?��B*��׾�̺uȴ��CA��o��B�Yl	��~��{0Q��.[�����y_7������(ߋӫ(y=E���Ų�"����b��K�����d�������HR��!�r�0��(g9r*&��`e�0�O�!M΁����.^tF�K#����m��P6j3�2�bç:q�(�q�xg��m��r/0E(kT�N��\������+K��9H�����oO�IU;�gg�1~���x�A�����ʍW0���bYS��Y�%X�.��Y�Z /���~�U�� W>SD�m�(l:`�s����FC�{H��>X}L%��IfǞ�ա�`�_�_t�T�E��Y�׵�,�%�����>�4޴k�v�˷<h����>����ҋz�}�A^#�Wu�y��}l�/)�!}�L��w���s��[RH��K@i�E���X�1���J`��E��tO�:em|�
�Jw.�2第֤�I�F���7�">�*�-����+ �����Óm�k�c-��Q���E.�4ر��͕�]i	��D��q�e�ؑ�CML�����N���c%�@�ȫ�$��Dv�*��#�E;��'�0a������!�in�P� _�
�p �J��I)�~��|���ޥ=�)�Q�nN
\���x�Wd2s�_۳�c-�l�M����ފř�̹�Yr=�j�eߴxȖp<T1/:�����@�.�HZZ�ׇ:16�����R�z� D��|��ʔ�>kH�:ˬ�܏�X�$��h��Z}� ��(�;zN��ߕ-�b�U\��K�+�!�-�}_�o�g鸜���c(w6;CU��w;f(�xD[.�P�P��g��:ze���hO�b�n�6~"9�q"������H�GأM�d��x�_��eD��7^�e��B`%���ϳ'�Y{�6h��\��^.*���x���~l^�C��,
��3a_._]���e���$��x��O�6e�=�D�푾K�H��r��vb�/�0A+O�A���&C�1>��6�5����>�[ȝ��y79r�z�/}C-���AB;O�jt8O@�������WOM���^�c�-���\�lG�S���of4�
���]mF��p���>���LW&��w;�kvę��@�]`9U�IS")�v����T;���ѫ��/r��k�ʮ��.{2�iN1�	��.x�4sT�F	�^)�B���-�I��F��c�^Dcb�3k����~'�u�{�^�
^5&K�f��EJ��A!�JA�=���nċ�Y@�{�\7�0ߖ��zў��S�
*��j-�~Ӯ�1�k85�!�����吀_��I�K�����[�Z��V@���¾Ѹ5�Ďf�a�:����6��d,0���B$LD��C{g1Aޥ��TZi��Aa`w��^#��70w0�Y̭-�
�����^�Ϧ�E��,	�\�ˎ�ɟ�:{ԯ4 �����ݙ�UC�a��?��o̧�:���B��>x&G��V�Gm�o���_=�J:nX�?�-f#}|���ٻ��+�D�SրU�EJ4�@WLH��G�>(ud��^i�6e����{
���(��l1��ŀS��(�fM3|P7c!�_(aA9Dq��&�\�ލ��Z4�1�x��m�{�wNԏ�
���^ShK|��9�!ȅ���fR��g�3����V}��G�+��R�/�$.�P2&��kO�_ͽ�J4Vy��Q���z㠍i8�/u�T�f���j���� ̈́��ٵ�˾����գ�/M�J�	��V ��L�����E��TldCVl�
�����������&~u �4�W"7΃��G��.�
H��A�ȥ�<��P�S��?5b� 9���SN�K-d��Q��B��/	Y�����/���m
5�V�B�a�F`���-�)�o���/�T���{�0a���ֆ�	A\��HQy�;�T��2�D!$ehL�2\�Y����, ܊w��l�m���jIM���I\����FL��]vN޿[�r����Q��Z�K�οU�b�-�O)��uLHDƓԭ�,�2��,1�1�wv���&�n&,��m
��~���e�V���!�<F|���Ō�(�+d�T�	���U���!+��p<Yd�?2��ϯS�K�]p���4G��7����
�cf�T(���i��-��	
~��;�s!��8�(��h��@Q��oʔa#$�t�/���i��-1[�&%Fx/�5�Ms��!�q�Qm$k��LO�j��c���3��sy�?�qw0���3����S����LQ�[`���+E>\�A۴�a�F�B[] r�G�>א (0K����-;�%����wo\��Y=�����
��.x���S9���j�
܉�1�/½�����9�VU&'���nOpo�Ct��c�^�2�X�iN�%%����+rB��Vcg%Ţ���1����e�:�u�j����Q�$��� ę[�fw6Sl+H���������r�@8�b8�C4�.�!�)bP��T��!�2�oθ+�����Ԯ�����'D�%{	�����N��/c���Ny }B�8�'wݰ�O�;�����D�	�` �_����j̢6���IBNF7و���o)�Tn�n�|Ψ���Y�������>���f��u�e���ő��}A2���R݄���D����Z�`#� ��Ő1-��ϒS~�Wt߭�iR�5��Os��3���u&�7���M*GR۱�q6"�Q�R�9m�2�.t t���~�3ޞ8	��,�ӎF]�ȵ*�`���#���	} ����~LZΙ|һw6x0J���u�%�Ž}�J��t�D��'����S���]�Nd��\$]�� �>�9*���8�y�7'�K��V��²{ g��vhX��p���21�W�o
�<�ן<�B	�l2��,��fG�`���ܳ� ڞ�)M��(��}��Χ/��;1���'�����sڸ0�#GIf@��e]�l���	p���D*�߉g�8���˺�Sq~j0y��\_m����1c�`�f,��8�?�� 䄾>M,�1��PFҁ�X��d%��u5=���ϵw����̷媷�>Ӣ�G˿"�<K"���֦�L�k�ܫ6��|��4ӳt]�[�X��aX&#ۦE���xuĦnWm��D�8Ul� 6kG�9�!�C�w?T�����8V9�C��C����,:V�GK�N��p)g�vL<cOM�~�w@L���Rz�3�+a\od~pD)����ܑTmF��O+.�s�׬�xg��r�`�� �6�`f�E�;{qG��YW��ǕeW��l4�]-�I�7ہ·K�5un���3t�������Eq/#*4�w��F�9�ҭ���DH¶��l�}�u��k/^� �s�%|d��� %�Ä>�g��(��ӝ���|�L��JO �^�1S�)�)�f�اS�&��e�U]�K�'v��܁�{����]Pw'�7���Q��6�����Q��`v�b�e5���G��Y�#�[�\%��b��:U�(`���5hܿ��B���&�t�l'�8?2 �M����:��`��$�	Bbz�P���$t�S/.�kAm�~4�R9�F[7�l���i˓���oMLŲ�zG�5q��k�6�X�O�A~�Dpu��5��Jz~�<G8�9<�<����y��?�\y ��7�]Pȸ��{��r�=����+�C���~~9�Ltk� 9�bP�>�����(Τ���<$�޶xiي��	Hy��qV���f��� O����-5��	�S°e�űԴ<$���px_�I�P����~�aG��=\Ҕ �K�����Ǽ�n8�r�y�~�N�=C����Ά%]rE�4u���]2~)i2!��ŕ��״�-��,q&9��:<��>Tb�Q�-~�r��qâ>��ʄʇ�^�?�M��6؛lὍ�g2�q���Rc�,���:���R�ۧq�j�X��fA����
�-ZqD�E�/9� OD��#է�b��dHX���#M��շ��s@q��{ �%�A�z��Q
O��E��V��_�rc,p����"��B\�@r�F;:�s%�7��i����Ki����0'����B����D���bz-�e	�|�٩(�R�1�:��/��L��s����H����q��@�O�ga�$$;z�N�5��X��z%
�,v�n�swN�۾��EG�����"gqW�x���6�U]'=~Oߒ������75m	�$���	�5���S��i��nc�sxa�8l���a�����A�bs׏NO�L�p2��Ǘ������+�R�g>��ֹ�䩻����5�������>g�J�-�x���V�uWc�q�O-��Z/#6@�+ۘ��s�ms��Z�q+ZS}��.�e�j'FԮ엂���.����=ю�lo��lV�L>bܴ	7 ��X=K��;��,е]3�U��͊�T�4��M�P��
��E�6��[�q�n2T1zSN6 B���_��p���c^"0�vK�2��� �d#`��8��� �т�j����3�}���u�'�%�Tv�8,���&}����+��ɫD�{���C�����]ʇ���O��yȷ����؏l4��	D3V~�`��9�$�����y[9Fx����K-,9���v!����Lܩ�d������}����蒪�b�T$���Z&�ނja�U!��K�p�"��X�3[���jސ��Eq���wl�ٛ��"�!U��6t�������+7�"��A�1��E�h�sS�!Iע�.������i�H>�?����Y\�KxtV�_s��d�	��z�(��s"��UK��G�ڛy~8�ٙ�ϒ\�7}��u�X��
~�eqW?K����H��|@'�^�ˀ��\�)���t;\/�[����k\X%K��<n]}�&X��u1ʹ��D&A�Dn̢��L�+$(x�k8��j@Y�ޭ挩��<��^}1k�o�e�����DS��6�}z��3��+���&ʐC�2��+�D�� "�H�_����`�4�1n��B���x��6����}�yI��c]kI��/��:�jQ�S<�L����&��Fp7�l�k��d����Ӊ!�$>�m)�Ή{��1�XQ���d�M��\R�}���M���aW3��Ls@��xm�_<R��>��/a���]�_��=^T '1~�p4�f��c��V�fa�a:Ţ"j�?$ѓ��m&Z��	�{���K6�gBY�Q�d,dc�H�){�7�˘�s@�h��<��;9$W�oD5��y�� =Q,�y�o�?n����lȅ):�RXG�.E�arB�E������!�����|c� ��"� |ߊEfXUҊu/���F/(�qL@�d@��Y��Dz�?^��j����f�B-����	D�W� �->�(ݳ������{阥�[��:�M�{�l?�{�bϲ�1��e����؃ّ%Q��Q`tC�D>N|�mP-������3��V)�2E��1�+o]D>es�S��G�E�#l6��|¬���`ǃ�p=b���gԞ0p	8���oX�(��F��?�׹�hDc3�פ~�����n�v)7��)�F|W4s g�)���5����l���f��8�����n��az���NoHŮ�"r�/޿��i1��Z���8jtL�~q�hY���.���6�?�v/�Q1�OЎ��ӓ�Ɨ�]d��$!��|�_�{&�V��Q��9����ݚ��ŋ=�,�;)��~y���#~�/ܷ'�E2��5��s�#	��z0-
�qR����S�������Ύ�CN��RD�F��d�f�,��*E]��o���!�hڄ����:�}���&ժua�^��bI[��-�P�0PQ�z�h�kkF+B�O�.I9kB&���I�o�yL�x������*��{�	+�#Nt�K�H�Ha����uė���HÃ�=�)�c�S,w�*E3�NO�\�^i�,ra�)FFW��	1����V�����:��"��
Xnp���p��?U2�WΠ^N��rm�@���h��*�LMF�v�ڥ���%~ojE����ȱ���h�,&@� h�p��QF֡�wU�O�F���9�/�k1i �D]����ê�#���"�ǃ�ݍ�~f�����?"Byk%孮~���J4}�=m���ԆL�� ��
(�$'5O�Fhc"��9�W�V7�ԕ���qq�;����S~
)D�8)?��BBi�<&P\L����^��;8}E��`��b�kKQ<Vj1��3"f5���yM��O5Eg.�%�޾�1]\"L�BĢ�uE�	`�!9mO��^G���i��5��c ��i��7_Wy�R�. �a��rm�Z��
�(��yE��$�fnL+dQ_r��5�W�4\�� ���3��7�h����0��Ƅ���9�`�Q����T�c�6�ݦ�>a_b$�L�Oh����{9}

8`�fHE9DKX�n��ޕ�e���*��N�X�P�t�����x�F����JC��ି���_�/{]sU���Ys��:�G�z��i����%����wn(F7�t=�u���O���@z����8њ��#�7+2�%�YrnjZ��f�ί�C�h��i�+�@c�'���8U�9S�w�9B@p��#U�D�<�T�IJ���
`/�l�ء������	�ϐę���Ҋ!��dP<���&��$�׏5�Ppk�D>�^XS{8��M>d��c(�_�	v6�q��Qu����g���׾q^inl�����;��E����+� [ב
/*B���ߦ9t��\�͝����p�y�fQAm�$Xn��n���{�K��A_�o��l�?�K�5y6�z�S��N]�A��q���M4L<�\�s���#=�=?����K6�Ke��]��s�O�� �Q�Bt ͍R ~�v�v�e'��Q�7�ݧ�/��>g�V,����g_�3��0�;�{}Dk�ez\����kj���X��,ǐX��n��Z�����Oj{=cM��rU�wK~�� ^��y���̋����� �L"7D���˕Ӻ��U�0�)(e	</��=��By>�M�!�����NŎ<;y���FU���#ޭh�Rr��IQ�at�6�'��BM��Y,^�E{�*H;ڍ̜��CQ�L���O�-8��,o�L����$_s>|���)T�R����5�O�2������F�D��9��ŏ��kم�ժ�<� ��m��ȶ(T[����+���Ͷ�t�v
��d�I����\���r#�־�`���$T��8�BKKN���S�-�:Z,zB�"9�^���ʰ�aU�2� �ԏ'�����H	T����緃� �1[�zU�6��x+>�U�O�y`(YdP� x��?`~���U�aAbaL+�+_�	��_B��������^@�Q�~H��.�n+T�9UGӺܛg��������x1�_!��gi�(1~�P){X �}p*�o.Ut���;ʡ�B�ZE�9��c'p%�et3~s=V�٭�g�8��Ɗ�PQ����_D��*�k�m�k����]��ur��ԝg=�-���[����^���0���+��k�hE�lg)<y�'�`���K3! �:�@�z&�m8�h�w����^K�UYW��V�qd�JF	��Ntگ���5����g	��;�疆F��tF&~�Q35�N�5��k���q������>a�BQ�� (<[�9�Ɏ�ºjk3�k�3B4_������H$��j�B2����"Ca=s��Ǹn��]�qm0-0�;���j㛋\fĽ� ���2�ᚑ��Rf���"h����xu��tr�u~%I�/�È�ZQz�Ţ�VM���>�/_
��UO�󄀰�x���k&9�G�h��F8��22�9_���<���>������V_X�G��Q(��9q�n)x��Z�5������	�2LO��?+$��+X;���E�CQ�>��]J�	R�����	�/�`�B��tQ��E��&zW��@3�uħ<Hw�XM4����v?Z�^	J��o���f!X�q3�g�ѯE�$Oɹ]���Ֆn�M�A*�Cp1nI$w�9��q�$w�g\�5J{��_����r_a��ǈ����ITE���[�}��`$�nB�Ϡ� �C��m|I�I��^�����׃�˩ML*�`�g1����g{6�j87Pc�;��Xհ��/�d�D{wN�F��aSHd���`Q�n6-���(�$ъ��GK)C֍t1��y�O�_�����d$S �����ze��������ֈ()�okߌ�r�".!�}ծR�X��q��&d���)������0��-����Q3(R�]�E�WT&S��ؠ����Hͺ.�����~��	A���J������'��^�]�c��W�ɞlW���E���&zE5\(�)�[��$I�`�Z=+,���<7B��g���H��[&33.�sK4�l�Ku�7Vi���N	e_;��{��q��g�#��'@Ϲ�c��h�
�Y� Q]�P�R��i)��}{d��|?��$QQ�2�k��;"�~އE��1�PQ�\� ��ȝ�-&�_������#��I�	G�N�(tէx��Z�-����`�m����[����l�㒆�������Fʎ����R��A�9�*�R����ڧ�c��-m�ȷp�h)ܢz}��Z��WwL�l5p�״�g�l���kw%��fk��ª|fmi~�QQ��RP0��H�'�.�aQ&�!��w6v@�����P�mI?�	Tؿ�z3����.�Es�5?�qݱL��>FC�.K�SL��J�3Ԩ_��Ԫ(H�f�J�T��8"]�J�?Q�v,1XH��o3��3�Q����������J=e�]E;�t�_|��3����ҕ8ۚG&DN�OO=EG���Ur
���S���H�=�:��u���d�֫7v�����ƚ�4��=�?�h����HV})�Md���#$h������k�C)�d.%���$����?�@�m��|�6s6�>ER���OJ�_�/�X��Z��A����r�/���ڃh����R��x�>pY#��^A��cO�˾�C)+y߶���_��n�q�ށ�(�0��i�D3�g�ل�RM��\���P[�[5H�[5M�c~�t8��S!����o+,,����QFY����J8)4�.͂�.�Y�����:O����xkx��Qs9��6��?�^�=ѝv����#tVn��S+�,oT.�K,Z�ј�TC��*d�[��C��4���O�+��
n�M�N.�7��	�8\��,&³�dCf9Ƕ�T5�f�0��{7V��p!�.\�I���/Ev��A�[��؏�.�ƥq���k��G��N�w���0Di�qQ+;{�t���wJ�o�ȦNu�o�}�`gϋ3R���O,K�Ó�X�� ·�2�����o����MH3{����*\�z4_x�&i����U����Y�GR�����}��[�_2��p�-'�b- 1�\Mp�H8������h9,UT���H[�b�|���]Y��e�x�#|L���?=K���v˾u�2���1C��1(��B���c��.�@�?U37tg�ƹ(B��\f�q��$�nVG�XH$w9fS��$jl�U�DR��׊�[����jK�cG��퍕�&H@6H�t'[��a�}��XG��F�'֯Ш���,W����](�a���}���/M���~���2@��jT��`������R�N@�����)���r�ʇ��0�`�p��qJv��_��`���P[�w�%���L�M���U�V��֟h�Y��#��e� �~���~:Z.oW�@9�PI�|ȔCV(�BJߡ���Q�-<ndaa�?RJr�� ���ŉr'{Â�64ƙ%aBO�ܠ��q���},��4Ԍ��24�mH�_���6?�>�R�ߟ��=nB�ЌfZ��BAˈ���s�;�������F��E!�ĐKRt3�!�Y��n�+c��{b�s�+P�^�'�)!K�Q.���F�0���7t_n�olV�C�95�x>-5�܉j��y�oL։� ��-UP�B�u7��H�ah8(�6��y��V�|n�0i���Lwa�C�Խ�$��#Sz������������/�ٷ�YF����<�����n�m�"���a����^g�a!g�s����<� ��1|ri�����e�����3��F�׊=���@��u�"��/�N��T]�����Zn��w�:�4�R{�p��W��p+��0�\C�a�k��#���ܴ�f�?=�������6�u4]�7�!Ğ�Mv��ī�����F1_?M��1��4#����N��z�hW��Kn���8h�l���Ǳl+qzVzI�Y��=�����X���P�� :���-���޳��d�+7�b:��=o�)5NQ;A��s 35W��v��K�ubFj�C9kX�2<�]n�#k���Sp�P�´���d�Z���gN�v!v�P7��s��þ���	����%xNAt���zG�ٗzC��Q�;%�|댳�`ωm))�QVl��Ņ��猤�j	x;��(���JA�L��Ф0�$[-�������#6U>�u�$t�@��:(�P�b��M��,��/�Y�6꩚Li*AƠ�j�{́�,z��(����(�U>�4���½T4�\�]�� �\Qpe}���7�y�v�����+�����B��Ǫ�޿�	����>.z[���N���a��C��������S�6@�Ň���KQ1�>�����+�����0䛦wbT{�/�poxQ�?���)?�]�N-�G��l��wN;C&���1�}�/�~Q�ie(�������)�ݼ�E�,�v�L|�N�N"�'ZԐ��� ��\G�TZ�����	�6Gz��7��� �+�v���Z�elY5�y�iġg����a]Y Cxn����>4�+�O��Ƚ�
+D�/�C������/b��Ѹ�Mb�l,�Dh?x�V��J ���,�+�Y�ь.S�*K�]� %���9��$�e�C\�=$���n�vC���L�^s�jHU�a���YU�7��t8�y�/eU����h����X�����5�ȧ�q�>�4�M���M���V���n�W��"�4�r��/᡻�,ȂFL�@nn'8�]L�1�s�Vo��FLj� �~�U,5�Z��9x��t�\E߳��rDPf�Š]KI&+�=�_ľ�4�U���ξ��W��Hr�岷�EC�{����k�%~`VoF1Fkeu�G4A�9��@V�Z:�hQi�4*w5�S�K	��L�R��]��v�Dr�v̾�v���z�Hxo�Ȯ�·{\�Qs������0i�MQ���Vo[[V���6A\��`�|Q.6���'Nx<C^\NH�QN�a��O�1%�^����.�޿���E�!�nY��m�w�$Qa~)Q�m,�#��Y�5��O5�C���菺�� �wd�P��Jg}M���5?�L�S]��W�)]xѫ�̸�av�:��@^����Y����K�k��
��&�J~�@�B�N��ųK1�Q.F{��c2F �	ؐf�N�*�!A��]��?L�鮋����Tn|k�e,���{��]܂���5c�!pBmd�5귁�U���-��$�~��shڄ� �.�%��U��lA����뚭��,�$Jp��������=��X�{R!�`��Ε�T!�`)�u�_�����-�,�e���I`sɜ��VӋ<��.e�9���� FD?p�{11�y�N����PU��lb�GZ��08q�|^קh~aǧNp���H˿�{�w�4��8�~M��vHwj���:/�}!���d���_c+����^l�sD�t|A(��u&���a+�z�]��2�eAЧ�x����"�N&�A-�Iuҏ�����%>H)��5��m;X�L��qj"c�k���c��!r&5(P�]��!�L��������V��^9��mxY���gT^HN�H0@F_�������v��ZAx�|8
�hit���d��'�4E�Q<5���b���b���S8eq[�iNj*�#;H$)Iq� `�l5�b������J�{���;�~_^��Cm���zd�5�����psC� fsqv��222yq�V�����uP�d�b��y�a_�me�a�\,;�T�.ƅ�,4{&��A�}s��0�0�Q)�-���t���ʇ�b�O7��Y���K	�-쵿������A�S|C{�Z���Y���U�2L-�'�؅���^]�Y��:�(#3�`'�b��6��y��7�Ĺ�\��tP����>[d�㛞�	�bg����/�'6����:���HE@}����؛���E8�(�&�q�lH>X3b�/�ߪ�ʱ�f!H[�uʽy܍!�#�j�k��*
�?�W�Pk>����� -��Ǭ�X�#C%I[%��������(�#r�fvi��Be����B�weTDa2�pr�����E�'T	�3 &�Je��Ja�N�e��p�e{�a�gi� ���� RKq%�H�K:��*	��U�3�#	r%r1��}ڣ�?��s���'L����K���]TXu��o�(�L�R�V����i����jݩ$q��SCQ.\c�P�C�{C:|�e����چ�VN�1s�fdqc߄D��¸��	�z�#z��02^&U(�)H�Jo1W��\1+�8�W}��P\��9�a�x���n����5��w�)����r��c��󾦌�<x�:+L���J��?ɗ�=�t�@�8�zGr�%�rB���w8m�����L^9���aC6�yl�`���p w5����?��'Oo�=��H�����u����IT�Sf��UkN��N��. ��l��Z�E�;���Y�-�Z�����&���%���&.�%��*�l0Ԓ���!?�Ғ��WA�xUA�2V]f�.�F,L�û�4��3�O�6&�aڥM~\'��sq_J杳��3B��&�QpS�d*�9u�n"�:@ڽ*v~��p�;���4gY�Y��A���΅� ���-U�B��u���Ǎ!��"ͦ��i�H\\��!Nu�fs���7o���f׹�1)��IϚ���~i'��C?{�#��f��k�Q}��
P���r)[D�b�Ո��E�4���+1!J`&��p�+K�l�U��K6��q9��^\��.�_��E��׀0[F]�����|��}���`4{�'�#2i)�m~XKAt�̵�B{:�J���ޣ�
&��C��U\e���������J������FD���jI8&1L�j(Gv�Q,�Xp �Y�.��:/�+�%��{��g/�xaT����Z����\x��4�v��!$8�e���s��Pq��԰�(����̸`!�ROņ ԂwIi���?�����W[�B������k�����v&��D'&�����.P� ��D�;Om��խ
�����7j_X��r�pۏ������_�6^@��95>@C�E�t}Z.��D��4�^.,71�ٵ�Ì�߀c���K�S�*���Wh�t^��ƴ)Y�sƼA���$�qd9cLr<*ּ�3�z�פZcT
�m�P�Z�#1sY�I�B3ױN��ȣ��)��Pq�(��+�6ųh������|9������@N�6Sm�I�b�
!{|.���k����δ�H�J�������^��I(���$T�{�/,#�5��ww��G�v�X�?������Y�\C{O�ނфn�Y
]�����ނb@=p�"��,>���b9�E٭������׆�
���v����l�xPK�.~��q߽��˘��j�YZG�ݨ���'�d�1��Z|�d�<dbs���2Ȥ���V��0��� ��caL�뮙���v1����|-��WU�(w�a5��|K��@�2�E���Z����Dt��3:��j��"��� �!����XbN�	+J�Z#����2��N�l�
x^=�l����GJP^&"ٓ*��!�*�m�CD��Yp����PR\
x{`w{K�!I9tl�?_���,�4O�l�Ǻ�����Q�Ǣ�}��Tu���\�6c'ʼM�(P��qF3&�M�Fiص���7�~�YTb	�jcݞZ��N=f��Wu����+-SU��x�2r�G��Q,�m��,)��H��D�����@6F��7�ŧ!�kKz��ݵ� �r�$����AoŁCW'i�hHl�����p����!����tBǫ'򀺥}A���@��* Nf��`M˨y8�q�?�����2Qh_�Dĳ�~�+-��l���i���e^���M A{rI�$����c6sZ>)��%�T
_�`|L���A���Z����0?�u��pځo%'e���J�ţGIp�(E�dS��1�7��TN��gm��H.f�)ɤ,�����-�{�%'2�P;�v������<S��/5���
���2r����������="j7~�5�qb��!@X[��u�[�:�:�
h��C�@^"�|�-��j3��I��c�)$���ISԈ$]�JS�3!��}�̆� ��F������x\C)�z�}0QF���K�D�XK]N�Eܞ�/uw>闕���-��o����}E�*Q���h��Y����AM����sp ����xYv=�Z�x��oZ���< �޴U�Q|��d��Eܖn�o�d��*o[�5x����T�ޘtE�,�׳a��9�'+��9���M���B滾�%	�bϖ��Ʊ��oXo�^v��?:��5a�w��K���=�8�~�Ha������d*����$.h��Q�����ֲ�LBF(�Amg��{]-"����MN�]��MBk׼�0xZ���٬((.<���gTy�;4�_i�.߀'�i9�At?R��D�}0Eg1��H@so��=h���M���~n���1`DK��D�Z%���B�~�:%}4���nz���#�*���vQ���^�x3*A�Fts�U�u����No9(+�K��q����g-���[��A�H��<~8������*1�Q�.>Yj����<5�;�z��<��@c�m\��Ul��a���8���1z0t+�ODpk���%gJܩOzA���!f_Ŷ���~�X�	��7�T8x1ݑHU�r�Q�����E�qp�-/�^�H|a�>�Y΂P�A�bqǥ��y%��W��m����aw�2�q��(��Xl�I+?� �������o�Ћ��e	�Q�m��=�J��ǰ�J
?�MeH��eu�����Q�c�S,D1�� ���і����y�1���V����&,
��������u��ġ�,��dm�Uk ����0��ev��U(���y#�0-�w=�4 _�D�@��>�Z��i8v���TMisY#zv;�?�~�[Ց١��^Յ��g����g�1^����~$��yG���u�H,��.E����>b_Y4�ou��k���n�FM��7���n&s��1J������`w��%��
L;�k��2S��в�}���Ty�U���(��x��تeh3`�u��W�k��e�ѿv=LJ��dpE�b���o��?=��WAGo��Co -��H������[ [�rg���6o��������.�ڵD���z��:�}���\v�*��v� �B֜�t�d��Z�=q��I����g�������Js�q�nf�n���Y�ؖia_��F@�V��8U{���b��aj \��lGM��|P9-�W*�X�����~�RY�Ҥrf\�j�bSU7�7A��8u�7h�y���d\��%9�6h�;|r��56;�,(<h�Ǫ=S&6�����+��B�+^K�I;�#��K��54�B��r�`w��x�fX�*��feg~7�b��c1���D4�g�z�G�-ԥ^�| �����%�'Ü@��1��P�'w���d�B�%� !��'�r�8`g0]
����O(< o�7<&(��zFLS�,h�Wo�T�5�p�o���rb�-j�< H���z���� ���Qv=r���`������b~�Y���A����I2"�XR��������.Jm�����(��|���X:Ȟ�al���Y�Ĉk`c�$��S�⫔����t����,�a8N���*&5��rO�Wod�Ѣ�,1)�%����R��OlU�Qc��	0Z�S�8Y�>���٩��@�+
�ei�ң�r���ԫ��ș:��}��Qq'�U��#��p�WVTT�L��&"L��Xe��S�ZG�P���K���u�z߉o6�������/
�������b�{�<����4�P�(�b��{�\�Ч���=��T6bBX�y�S�y0�,�*�]<�<
!�Qm�@��P\��p4굎PDF���g����15),�k�P��U������Qc��]��,a�_���%���we�����I�00�8�Z	~��u����@���V�/0�YF�D��	��y��޹w�&
꽉��M/e&���+�@{����g���$�K����eV����"����b�}>�0r���M\I#�d+����E���^RC}�Rz�wٖƨ�p\k��m0S�.���
Y�/j�c�cҨ.�]���m��սto}Ì@l��ǲ
�+�)�W`ɏLУm�xm�W��
�
�w3���2#X]�,��9�+�,�U��*¬�"p�,Am�x��l��w?�T|p��3�mL
�iD�j���=��x��d-n�����
��*GJ��}�#Ӛ�;TV����H~��Sao������t{8zE*&:쎶�:��%�r�D��X���h(f|�v��$�U��Z�{o����|��DY[�f��fB��ǖL�������S�5P��:	h��D�4�'���.�-�z�:1cg�>y��Q���h�A�ɧo�ѠZ��$+�5�,/���o�^��)9:N�C�q?qӕSk~�n�l]ܱ�0'�n5N>3��-ٔ�����B�G��1�p̭5��ߘ��|͈�._܂&�i�I@�����L^u����r��Bd�A�$�I�ѡ�	�}���sPrL�J����m�
��d�^�"��a���A�5��9���q8��&��ֿU ��� ���=�2%[��68v{��\���bP���\Ɯ0B���^�z�S�ǵ�hg|]j��y��(�n{G�$���������ڕ��-�1#����NM�������� ʙ�eVQyo��0t���I�a׬W��`�丗_�����5���@2�Y�gg�g��s������zY��4R5f�� ���9�c�=�?���P΁֢��57�T��%�f>�r��9�+�����(Z�s/����K�4P��\�`��O�$n�\�g7�C���2��.ʦ#��L-e]kº�e�)b��-�#�T-����/��o�$+o �A�=�r�]
,$M��Kg�Gt�`����?"KL+"L�a1�̋����|�u��-��A�t�4�tO�(�w�����9��S�8{Lۉ6/��
ԛhE<�!�i���9u@k��y�A�����^?ZH�]�

vل���'�r��J(�vN�E�Xs!���]�v�U��>h%��"�p:���w5�2��\�hӅYR~���\���2���U�������7	 �İ����%���g��b���K�wӄ�h�Zp{ ���?�9}u�R�^`�h���[��*���&B]��zѶ;
-�~x}hO�M�C��|��j+iAy/�2��o�%zot��	nq(a�Lܲu�lF�~�oJ��!g�k8}N3��-�Q"���LV����O7X�dSHb`�G��)�dW]mY�kt��X[Ȳ���O�.A��{p{��ǧ�֓Z|А����VеQ�A���Y����w�M��;�I)����Gy�~&��^zh���#��k��q��P�0�G�T��1��g�KDU26E��b��H�����!ҝ1�B��d�JgGhm�i��v�t��ҾW�����j�NĸT�.������}+h�T��2���ǎp0��է�F�n�i���KN&=�"=�=n�Ť�z�J��}��~��,1ͪ��'w{sg�u�ʇ�ǻu�0�-�(G�(�Sa�.�2��/UT�՛������H��o�G�ڜ�Mĕ'��F6Kځ����)ki�z܊��o��QH�r��M�i�����ZX�@=�(ж�,�擌�L�͏&%ϥ����<���wnO�2+(���&���ܑH2�%K�J
� ^cJ*&�V�P�������t�t .j��w�`l�eΟlຫb�;�,+.ʺlk��� ���Ӎ/� ���2�Ϊ���,)�<�]�c� 7�-�m2U@� C`�r��3����-�1�(�
�î﫠,�������hiX�u�����3zH~>F0�|�p�X����q�j�ɮ��$��f��)��/��p�Z^�5��r�����/fɨm9�覟��5us��H��]�X�4QZ:�w`� ]Va7��F�|Ҟ.�̫���	�i�w�R�S�f��Q1��l�[���".~K�Y�������HÛ/a�"��8�7����١"�j^ahb΄ߠ�W�=D�Dl�F���@,�����%1�#�G�d����-�Ͽ{�h&F�!��Ҏ敬�bK�ϑյ;YXC��"S;���V����v�t}���KW�J�2Ý{`���0�`U60��K����(�`���k�=`�6���d��4q�'�F^�s(X~����M2=��$�g�~��k��k�,���B��՟@VG�P���I�)��� ��̸�1^���)��bck�6��I&Y�.�'��I�6�H�t?V��%�W���C��i��&mLO7ٖ���`X`�ǽ��$ܨ]�E�F����J�?P*�r7�����n�}��']�v�X��;{�"WC��Z��AD�%?NW��`*�&�~X���'���n��������S���o9�ޢ�L�2����m�铦7�B�������
��Z��7ޢ��9Z���4������%!N�O�3���R��/@#L!V ���\6W1�`�if�/J�yT�Y�QF����F����˟H�6N���a١.$1![�$5n�Z�yР�eE��6y��%�h��ϕ���uu,�������|�!j�l�������hR���4�dY�C�ؚ���ci�>i�OW^-icPF�Ѣz҅��`�-1Zw]��YH��22��d�B./>*�=�d�,h�ێp�o�F���*��?�|�B?�;�6�]�� e!O.ń���Ԑr��_w�B�����4�Ct�:���.�ӎ�60�dV�`�u���b%�J��A�������4�m��!$gpu�1-ld���Vt)Ǜ.���L��Cr�c����>�-�2Sր�f�|���`�B�)*�8�?�"hL�B�ùU��|�Ӄf�|��/��PN�WV���%���d~�f?���<��<�����Ŏ��c��̊�,J�ƹ0M�
�H��?�
��Ɨ߷2�r��OYؖ��^A5��B�������ɟx�E�y�*ۓH����&�4w��Z�VR�X�b�$V�g|��ř���H�]�S���*���9�(W|T�"��j�jD�>���sݙo�b��\��qz:�,�)MУ-���.5	|E��fC	��C�ci�UQ6�n}���ϳG����{S��x:)ε�������
���֧�Z�^�JX���2I�/�V�g�{#r�2(	�]وE� E>�!MS�X�[lh��3�.��qk�uD�&��Q!�?48�Sn����ѓȂ(�]�|�2�Y;L����56���ˎ4����n��z�Ƣ���)?	����DSd�$g�Ԫ�;滟�ȧ���r*�3��o�|��ZI���z���ک�<u��)�D��C��pJrt�!ǀNj4�zV��de����Z�D�N
��P$����x��`&���ud���[3.=w.	w�͘�2z�hX���6�"��@5��o^<�@���K������f��жl��_'A?O�3XIi��4\G��[v���8M^o�G<���������#�ߗ-FZ'��D" ֽZI`9�1ڗ����d���E��'z�7�����_�E/��+�d�u��]I-j��0��W�A��0��#2�\B�Dp��;  �`�f�HF�=lv�Ų�����g����y��Pw|�.W��'�6v!�>�D]���}$*��5$�@�UDY\��]��� �� ' M�f�=> jZX����Si�"lr���m������������٦c��kk��m���.&Ib3=U�V0º�Ê��6��X��I �sь/
��m�AY��W!��Z�Atb�θ7~"�t�8}� ���0�&yoΣ�ȱq̱���.1���mxj��	Ň�4*��%�[�Y���\.P�,\B�֠���-zo��|8|:(6p��Y����<�����x9��3b;��	M��ѻ2��K����'׌A'�&��1S�V��wf�d���+O9"��R�]��Cb�p���/�? Q���|�����7�_Y�1��P(�^�j��yҷ���Ѫ��k�)��uq�g��bJd�;������c����ؐ��6P��g� <ا7��k���m��g�����ëh��F�}�ūu�
@D7�g�l��P����7�]%1�L�2�\cW�H�;޽�e�J�Y��:�Y���DđΧ�(���㥄�&��!4hu�H֨ytF��+H_qf�v����:ҕ���4�O0�AM����b���>�@U�Pb�ϙ�{���r�2�����(����1��<�|4 |����5�N;�/ ����M�����D,AζI�[o'7m���W�}>-��1�֓��Q��vpYj!E�Fl���#.��|qRH��d̈��rF��0?�n�b��ge��-�=8�@BMB�7=�n�(�VoT� ��(=fJ�z��? Sc�O�ښ̍�ND%�����[-�n�Y}n�:Q�;�)5���>%hK!�$�b+�Z
n��3��aV��Jh|�����I�-��(Mf�P�E!��
����p5�-_a�`�q+� �E#T�ؿ�.�:DS�� ��_�^\�Z�l
8����g�x�ްc��&�g��"}L�"�����ɽ�yUq�Ib�̛��G�C��S����[�?޹����2��<|f����y玵Zn�r���8��co��YRlj`�с�ٛð0:86��L�D��Nqp�F	ֿ���ܖWn-7��u�H�	aZ�e�\�a������ؔ W�s�/��|�i����"��Z���Tls��->� )�+��p9N����E^lA$�����%@�߱����>�A$����}����x^z�ҭB��h�Z30*F��kE����z�iq�eG����1�w����I�J|����|�g"�Ɯjf���8Nݣ����͒g�
��H�J[o ��D}d�U� 3��l�E  �Nu�4�V�/y�5ω�}��0��G�:�*��'Rzy���K_�Mz�#_.�9�B���s����/淊�OӅ9;��AJ��D�ė�=��6J�V����٥�1<n,A}�y8�.�kMA~nn	k:�qPj�DI�����IwQ�uFʗʩ;BՓ&$���� 2��o`���`V{��)q��n����Z}�벸"b���Z|�D=^
'x���|F�8;y^��Ҏ�ߴ���~�]z������	�]�;Ѧ�2�sNc����[۷	Z�`�?�	9�/�$�"e���=��]�^?���=w��	�8|| ?��ISغ��"a��������A|y�c�MwH��pޞ�?���c߇�y���斀dx�����5���&���`�.L��Ш;Y1'6���ԯh�<�����vN
���]&�!B�1�@��	���,c%?X$<��Ī�l
�����OV!���ّ(�05aB�+�3:���g3�$�����2���W(^2 k��.q �^|�Sh���u��Ӫ�t� ]M6e�&�eFy�AxV>�&a���@�?���X��u��Hi�a�=�/գ^ݹ��/�F$H~��F�5w ��/�/���m�~� =P��<���a���	��'ؐ��g��kF`��=�I�6U� e͚Nh;03��3��Ǩ)!�ɀC��R��3"��vד3�#C�z��FC&+1����So�*�4�<}�� Lb#T�o5P��P�*�aVƗ���B��?.��U�H��ט_�No�D��M��:Ku�;������y��@N�y�==�*�K�,��w���-L�>x�&UU �'��_Q7����Zg�ºXG��*��P��*�XG��@�\�r�h#:�1�1��xZH�F��[��$��HW��6�Ս�수*az`*\@�	a��^�Sr�ܱа�.T�4!ڹE�,S�{��}���R#D"�/���I�2.T#��Tk�=
��j��s<s�|���>������M�<�é���K��[�X�ն�����օ�h��X 1e_Φ\f�x[hc-�]��cm�L������� ��HmXLur� N���.�-� ����<�q'�����\c���W�t1�4)�Х!��fZ*Y�\qt���[�s�mV#�aE��Z���?M:-Ӝ�Bkh۔�̆&�//:��}��cHڅ��ޓ��phA�|,vL7�T/�Ω�_ܧ(�+t0C]B�)�uT49n�Ӄ���������Ke���ANT�A�4����z6\�
Q��HĒ�<~QK{�{��/c��ܠj� ���pz��o�m{���VO�Ya��jF���QH'��6{)Ax�m(I�һ�2��D�N�f-M��ݧ�Ǟ����c��2/���'BםY�h=U�~H��#yRm���|��h.@ăc>Ru�ɇ�:�ҩ��_��n�T��˟R	�Is���{(>,f�0L���nL�R�z�����f�����!��0�8B؉\�!\�U�o��,`l?���l>�i��E�;�{��Sg��/fL�9W�!;�J��#����8{j���ߵ�Kݎ5 ����(`){��='��0�hjdLjR9J�A?��p�J�"�.Z+�z���X��^Ы��&ԥ�O�����K�����{���]�[�����>�����[�zgv��kc�S��-9G!�4���W1�r}�e��c���P�����%B�C��V�Ԕ��'$-��i7(^��CU�P?+I�W�"��[]�P��r~�,=��)Ա��U�5$B��/�i��'�tr���4�e��,�,HE���q����D<��D��[�0�����������r��R���M�κ�]Źp[�*�_��ǝ`H�С�'�Cx��)��T�~�M%�FfU�e]G��pd7�����P3��W��8�@C}�8��Zm�4�d�pUp�aԦ13�)ӱf|�1�˿r#�*m퇫�@'�#���Qr�+���ǚ���p_�+}��Y�b=/�=�jH]V |a�3z1�P(�K0���n�rg�
K�ES^\buj����,��>&� �-��Y�qV�d�:m�/�	���gL�I�I߹u����jڀ�cR$'
L�nA��o�W��m刃�{V^Y~k����4����AB<^t%%���"�7�<PD�e����!\M�K_Ԓh��΄-J^��#5�iy����`�����'��4�[�T��TT�j-6��*��s:
36���b����P�N�7^B*��x!��6H�c�l��Qegw����Ue�:�r��?[V$߄1�m�@��'�e��)P���E�e��*K|�9^��1;r�g&c���I�-<ǯ��b�ՌK�����d�����*�^�w��\/�8�ґkɆ��nu��Ť�R�a���~��9��\[ͻ���BPҦ��2��Ťa����f���I�	�⣙=�Ɯ�{��eV)	܃hRj�\w����Ks���ؤ(��b��&��w��x���Ϋr^s���XH�Dq��͌tW�a>��z��Ɗ��#��f�t��T&>�\45:��d�X�")�Y�WAS�a���w���}�t����VC��fp����IjX��<w�k�`!Ш����sK0UC��1�����d/ar�#V�F�����垄�Q��ȵf��p0�-��Q%TT�f�*��S���a��I ���3ѵn`MC?�*Q����SS����ܕ�*-�c��:C�j�.CvFI~ob�}x�Ɣ�C���&��'���@��%@���ׄ��� 6�n��V	c��e%��s_���	^b3O������2�&��$�����S������f475�]3���f���u����j��'�t�^�de")_V<!td��̣8���B�zd�O�u��(���w�B3��t�%]�����n��u:�����_�	P����Țs�ݠ��+8�閖{�F��-��uL�'u!��FT���)))8��-c<��}�T���Qg+�C�R�A�j��>��u��U-�|�:�*NU"���r�&n�ꌅ������.[m8I6g綸�o��H�+�kZ҈
qH�IO�ef�)����Q��KOn��Y�|�5�H�/ai���l����#}g��jW���Em�r�9���X��od'�� h�/!}X/JȾ,��:�*{�b:\�Lk!f���N�%3�.�N�VX�ė���O��?з�!F�$&�a�ׅ�@;�C]{޺�t�bd�:r:P"�.�p.n�Rf��/�
 ��27���kX}��ŏ��'�&��D����!����(�}�T�}!tȬ��q��4{G�>@�ĳ�'�F�C�U`���4�,��.����6=�$?�
]m3���;)I��]��n��H��D�o@Z�+7��w���lb7���T yj��v](���¢h�Ygv^U�4��)����m�V�.LZ�	l����/�@~��tGZ(�K�Ã�-f{X�mW	�GM%����?��ȃbWb	�n�f]�8 ���5(�����7'�L���'g���F�47�xt�F�l�s��g��_��h����6���-��|�:3��fk�ֱl�n�*i��uK��|FC͒wB�<�H5��V#�*��]8l.tg>�s}���y����Pj̍�<m����G�\�oF�m� �;P}�L�,���R�g�X(�{��\@�m+Z�������[���G43����T]c28�ˋ:v��S���+�,	c~(����{(�.xw{�7}G9��z����j�G�zy�O=�rf��o3�i����8�Z�1Z#�s�&I�c���R��S���Y� �zN�*�ߟ�˕\'����i�{��yڰef��!�o�w�$�

��i�,*$�=�R�?�����/���w�@<��q_����M��6u9�`"
��eȥ���[���@T�VTR�!2!�g+��\�߾�m��x�zV~��18@��خGfD��j�����B��ڲ�O�Z�V��ܤo����5S�����3J� L����w��i���M��#�5$�6���=��|;�[��MD�'�]�q���K�}an�a�4�t�E�}}���?n�e2�X�CL����r~C�`�H���mCt_SQ��*OZj$���f���6�wZ��T)[𕉴-���fb�; %z�`��`�,��A6��K�c<@$�'���T��}%�X� �(K�Ta�ӽl�X�U�7��X#����	�������9�#���v����!��Va�,��>�/^P `^'���,�:���rX��P�kV_����^ɬ(����<���1���!2��hZ�z�f�m����b�]��;#^��4�6���>r��Q��͉\���<�3Ǧ"ȕh������=�l;-��>�2��8)�����vn���-�G$C7PE/L�>�p�f(nNe�3�L<e�@�Qߖ���Y�e!��Ң"B�f��:�&�UfD6１l֗���V�����g��׵�u�n\�x%G�	�4���~�k�ʤ;�.���7��UkT��Ďz�x��_Y&�)�)Yw�d!O.��X� �	E��Z��=N<�S����_�#�Gߌ���~r?��iM�(A��)��	+�����r������f�=e�3X�׽N޿T�K4��Q�b�53'�u:��3�ٳ���oH��<S�i2*8�ja  BϹ�~	�������Ɠg���}L�Ac�1Q��Fch$r>�k��@���+s�0��4i�JO�{����M��WX͇Fq����m@�T/<��'��c�
ғzބ���j� @�;�y,����f�oloq$�/��ijn�m��k�{�L'̸��_|�=(��;�}߽��*�*�fX�R���3Z`]��i�l}�����!��~xi/�ۏ�^^�ks��	+�ht����ۇ��@���]���ݿ���M��d9c?���.g:q�A��Wj��#?;+�6̺�'�5_����I:6�b�J)��"�<��ȚH�4��Lag�^.��K{�vi�����#�x��G�� ��omakL{ }�E����s������7⁍<$X�ug^��g�A���CH%G�����L\���ȩ1����U�/^FPx���['���'	�L��pVi XiybU��<$)%C��]��H]�b�%��8�ن<�7ƹ+y�+ܘ��"	G�2+kc<2��Ucܾ�E�=R�1����_��n�X��}�	��)�ޜ Z�}�ߌ���9��΢������B�0�1��+G�g�~�5\�<a��*�H�t�RZ���zE������D���zç0�*�!���������b�	�
 ���w�j$8��i�%Й�δ3v7/�|�u��������@��hv�x\��q-^��#h�(��X,b5���aO]8UUu���鱙� ���Qٚu$HH�DІT
�nW:gA�i9��.�-�^�N�4��Ol�d�x�������0�]`Ӗ�T$��k�?�б4v�'w�t�/H�# �p�(�,�}fJ2}�W_]��.Ϻ�;|-�ݡ����v��k�6n�1_��+LK�ֶu���hK��{�r]�|�)Y��v���c�B+�4��Zѱv���X�/k�i��Oi}����3�`��H���vFX�bEl�=@��fw`������1�3���g��} ��h��h�'u|i���%K��|e�G�`u*%�"��.��&~Mh���rSϞ���*�h7f���$�A���%@��n��_�:HMߪ!��:�Y�j�ij��xts߮���b^Q���ˍ��0[[<�>Ȯ�������'�b�o�rg&dksw�X�0��KS�h��l�Z?��d�l#�S���6��� �<��c{Zy���&�g��W��c�MJ���;�M�v"��	���ɣ�����8⚥-ѧ����>�䖶2ᇯy0��l����H����;D�ֱ��뙪K�rCX�:6�ǋ����v"aL��М�~�I[EY����H�/�.r�c���++��,制��A���,�0*nZ��c����1q�}���qII���0p
�N?���@#u' $g��6�{G����� �?{(���dAu��/ˈИ�q�q!N�9���C�6/��'���R�����l+�Y9�6���ft4��O��j��͞���x��|��� ��@@��u��_�Rԯ�-�BX�o��2u���t�|�	'0'�n���#�W��Wͥ�cc����Ԃ~Ǽ"��H.����'}Km@��{��D$��[��
!�=��P�s��r�k�)��H>:��S��(��њ�޶����^���OݣJ���G�bA�ǘ%'�	�(J�[�d>��=v��X���i7�Ե�ǟ* ]�v�A��*�^	az?�·�bw�]_��f�/�Us�|�S���-2J���w�#��
��gj��qᧈ=Z�ฐ�kb�<t'�=���"L,[t��^��.xސں�=��0�D�D��Ai�l{��gZ�k$�..��C�(;_�7έ�I�>v2�s�v��H�26�U��?�7iQ�ܱ�n���B���{�������M����g�˱�����q�4����ݹ�^���ӠL��(��jǱ��i`׋Y�%�B���P#��y����7�$������t�-(��T�GmvKc]��N3u���j�ڇ�L����b�EK���G��.R8I�rZ?��}7��f����������qX�2�T_�y��P��!����Υ�'�����n��p�&�W�J:��ru<1��K�Xr�0��R �{�!뼝v�"����ݢSW�A$�K��ll�6�����Kq�9ym9����مX�F���F��'���'^x��ڶ2=p�beA��MC1��C���;AJ�f6ަk�2%s�D-Oz?���<v���Ibw�V(����F�f��iy�^>�l�i��J��J�����h-�������W��F�8�(�Y��`�ER��q�e�����0�B��بg�����ېָ�ZIj�{8�s�4ت��f�ƒ6`TG1�WϿr�u&s�>�R/7Wֶn���
�'�M��`S��V-��pn>��܀dY�	Q R���nv�C����l�E)(��VDLn�AO˾�]�v���z4_>@�{��(?���J�kްل��Y��P�����$�G�]W��5* �>��CQ+�7��7�����3��\N��n,3�wFR�����ӈԴ�i�������Z��߼9�G��6v����{���������u1$�2jN-�K	��G�'<�ϴQ�����y���*���M��S&�����8��~7�!2nǰ�aS�h�8�Y\��Ѱ!qu$��ƫ��3��9��K�=�6���� �ĵP�3�!���1ޑ������H�ʔ�����!��!N�|�!"�nb��"��̿�]W״t;�#��_����;���:��g�תd��p3m���v$e�PHbq��1�3�S���4��^�z6'ы@���%%\�ȓ^%�::�`�6,aG�C��׊Y�a���hD�r�br�J2�BM{	�-��^ �>�Xi&ē=��"�S�Ti���/w���]���٧�V~;M�%U��t,��vwYu���`O��a���l}y냆�Q�XΡq&�w����'���8Ѵ�m[�fB��¸�-�1�`Z�E0�K5��֘4�Y�	�׶�9��C(G�j�~w�L���?t��TL���'��B�U-�r��O:Łȇl�����Ԣ.�
nU�o�8�&��[�����5!�u��K`Tk;�\���T-&?|ǒ��	�XAu��f�k�(=R%�ֻ@M��**��e�������'�����̤�W0�՛;(���n�^�z8^|�����zaxGQA\v<L<�/�I�o/���r�Y793��Y�o�*ߴ\�ʇs��ᧅ�?+(�Hx'�G�;��SC ��ٺA�K�ҤF��^,[l���g)��Q���+z�n�+�t3�Jٜ<�S������92i�b�7����f�WP<n�e
])(t��Z� ���A����c� �2�d��a��^�Mz$j�vn�J�")��W�ח�/�7�Ey�e_Mms��LБA��w^�όإNcq�c^��}6I2���{�<	���o�]?�/��C��[�qY�u�R�^�!�&^'�[��Z{;�dS�|�3�ƴt
	m��ܣp�B�	��`5}o���>�HXT�,j0јÀ�$��L�c�p[���h��j�w!�F�>�!�#�fzʙ�K�������qa��|�H�{���R�_�=Q_S�K r��+�W�`�ا��=������J����&JꘜMS�(. .ƺ�wyAȌR.���R�"��	��PK�ΖP��7Ƈb�n���oYd5��h���i�iW[�ڛ���[R-��vDP��l M��$Y6݊�i56ð~�	�4o[��k5����~����D�cYX���ϐ3wK��SԠ~]����2l���[E����?�f��C�\c�^��MS����		�~�v7�d[wcE�Z�-H����A���21�=��z����.��v �Ħ��ҏ��3�.�'H/����G��oDC?K?7,i����NSՅf_�;�1K�+6 ܱxlD�(h���������&O�e�Tm��_�S~� �F3�v���2_���T�ӪX�H�����ǹ�Y�d��ɺ�*���5]���j�W��9��r�^ıڅ����=��:cќ/�`,%z�xm�%_[e 0?ڙ�O��(�/�����ӌ�rx�u_Op��Ϛt<�Rd ��õh�����Q\�tf���U�gXl��ٵTȊ'j������S�:[��$��5�"�B+�#]���]����eڝ4*l?�{��|S�>"��"���E'w.��ˮ?����[)��,��z�И~+P�������pJe,P�^��͠�N���a�C��D�B�S������6:����i���{��""5#�b(����a��n3c��w�>&�r�9��hS�������%�_�-�A�b O�
ka*ʖ��l$��Sf�hM�Ç*
�1��muظ��M9��Pk\~��`�b�Rj�.S=��?�mM�C)ۮ�_��I����\qq�QcJ+��e��g�*�=hd/�VS��Q ��;��qI�@*��Վ@H(zX>%J���J&����&.��L�-�������n�,���;(�l��&#_kx���˧)�[w����VEyy7!uS����5��
�Bkp21@a�r�����6 ��]O�2��zO��i��Nu����F+�Fx�_����Z7�ш�-R����?�*A1-�F�2^u��e[MK�cv�s�����~gi魉�Ŕ(������wm��k�az=�i[�6�|����T:$I���@����Y2M��T{�����FFB�r��3᐀cM�1DE+�ꪬ�,uބ�Kf?��t�{�U6N�ڊ�I��i��Tp$΃��n��w,��L�l|_*v]8��"��_�� q�Y��,7zc���U,�K�|:���>�`��k�V̄(�u���z;"%DIt�ɑ��u���Q�x���zh+4Q�g���F���č��Qh��x�Z�:kf������+1��=�&hqxPvfHːy�g�� �,�n��7�c�8h7;��g�W�����x/�����'�7]�*Ȭ��0���/e7Ib���g���
�������vÎ�]�U�������w���Ƚy�F'e=
{B�*��ŏ!@M>��p��_��g�f�i��v��k�r|���Ld?��B7pu��y^BUBM>;�1�VUs��~��ևD��Oq�[���\�� �bt���)�}�,%QƁ�����L����OK�HB�$�2CDYk�����쥨�
�t�P�CLߋ�8�y5�Ib�E��Tz�6-WɄ�J������5Vp�>����E��D��Bi��v=|k��-�_��5���0��;M����b�pla�D(Z*���ѱ���6\�J���ci��΂��&W:b�_	`�M�������_�o���\tR��#\,�K���>�v�{;I'���Qrx�,������Vy�C�6	��r4���:Fd�>��]������?&+�y���Ֆ6�Պ6��n�Ġ7���6���BIk�X��	��|���|P�,��6�|��Rr�� �e�-l��^w:Y��"�uE��D�"��D�ED�|k�E��`8�0�g3���GY��M���p&�>R�� '_����Ɏ�8_V��(�����c��U2�G7/V]�����ڭ�W�C�����d������{B�zNߚA̺�J��^��{�N��'`ח}����}ÓʩsIh�����-i#����g�U�+��F�c�4U9�#���M�T(��S�Yi�r�tU�I�*��
�YYuY$N�"N�g�n���w����lH��c�)�1�$��R8l
~��L�l��b/�~���q=V�G-P"�	"��6��f�'Uk����r
%R.W��k�N�$���Čr�:���-)d�L!\F)ܱ�Ky�[�yp��!�?K�v���'L�sEI�ʁǇ����Q��>sv�O�:q�t��J�������7D���L�	R�D5^�T��̪swѷ9��b�a)x)_���|l������YO�w�	�ܜ�U�g�v]������7L����U\e:ͱ�����࿬|�S*;$�H1���Jڱ:"q�9��95�j��W0��:J����l���s��K����P қց����i"��Ă�n������D�{�.WPw���W�b]�>ߧ�Q�b��t������������+�Q�b�|���C�b�kfP��*�D�2�a�Y��*���Rk�3�Z��Ø�t�]��n�G@m�:	 &VU�k�;C"�=�o�	86�lv�yW���UGF�xN=��.t}�=iGnvrj��� �,gH�&��g��wv_f��������b�-��M:��M�.(@�*����K?l�gy�F4Qb���4��̃U��P�T���*��@�*	Sha)������&$М�7����/3D�� q{
L�[E]�<�s(4��5j�z �k+�Hm!>��
`���Qdy��r߳�b4Fϫ��&Y��K���_��,Beh���b���p9&l]b��:r���F�k�7*}���*��x��^9[f�+|���r�3��Gߩi/����YKK'ڐ�Q���w����_��M7_���CE���e��7J< u��\�Y��+[�e��\F��4A W��c��5�  ��ҙ3^�Ъn��s�o���b��7��spR©��p���µ���V�x��������
��Pn�yt�%�8g��� ;C}�?�&�{fȦ�S���^O�-�F�p�����䮣�-1!�{���-�䈰^8�Z�U;��l�;���q��� �E`���[Y��fy��\�@�~�y�9���7*�%�X�s$��w}��&j�-�g�8�;�!�PZ����[S�q/�4��BW8��Hi��"Z>�*A���Y"�+Nĝ���]	w�]�|t(�P~��A3��x/yVh#u	ԗ�?�9��8�c� ^�E�C��ʋMT�A��d)�#"eT+N<��r3�%+����_�<3o�t^kH$ߝ7��Ւ�;���� 	u;Bm@�DM
�U���D(�`N�jO��Rs�8��L�u*U�K��fq�D�]2�h���\���]�9M�w\]^�Ǜ�hN��$��CC�1j�Ќ��W���Uy\Bw��[b�3^
��$2�IO�C��;t ��E(�zf�I�	L��h{T���1��KOx4tI+8��/�H�`k*l؉;�Kc]���Y;UV�n"�e�o����9U�蚷��\�ļvY��}��)�����S�[�7)
��lg��]v��ak$>Lϊ��R��Q������Ϯ!�ԡ}#Se�8������7_ �~�I���3A(�쮄�^E�����$��X�f�Q��[�q�� �%�-��n�e�a_��e��C��:�Ed9���g��W2���+np`}ka\<����o���ף��T!Mqif���ۇ�loD����#�Y���(\X�Li61�p�)�C���,*�x�=������U�Y�X��+���7L�ˮ��=-J1%7��@	'�-]-(z����d-B��K	/oj�8�w�$���4D�NJꕀB?�q(�8oG./�F$r�fP~տ-�8E��MYܛ�_�����a߆ۭĄL�n^����	0�>��K����
~��z�����MEmW� �j�]�G����/��?!�:A��>9+KWKEָ��[���0X�Κ���%�v�l����4W�}�(�z{�<����z���^�ʣXH���]}�����^���v����oϥ�Dck�'3�1ژd�Z2�MB�*N�qc��3�X���w9܍jD|v_�Q�|��f\=�}�l����j���!��6��~yw�?Hގ�� |��O�`�ι�Mj�𭫟`�X��dx.-^�5E��ʃܱ����Z�^~�A�Ρ�.��q�_K���˅��J'A���U�3�w*ۀ�y���֡'7sU�R��;���u��l5E��`ʠC�|�P�𦫱��X\��S-O�(q��5��5���YD�rt:a
��a��2��>�ۗ�9�/h��:��i�:|�m��D����%�[�8��wNnS��&�}��������ܴL��bPz�c�.���O��.������j��c�Z�iI�����A��36@Y�lWRGnE